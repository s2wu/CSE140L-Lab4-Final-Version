// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Feb 28 2020 19:07:29

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__17566;
    wire N__17565;
    wire N__17564;
    wire N__17557;
    wire N__17556;
    wire N__17555;
    wire N__17548;
    wire N__17547;
    wire N__17546;
    wire N__17539;
    wire N__17538;
    wire N__17537;
    wire N__17530;
    wire N__17529;
    wire N__17528;
    wire N__17521;
    wire N__17520;
    wire N__17519;
    wire N__17512;
    wire N__17511;
    wire N__17510;
    wire N__17503;
    wire N__17502;
    wire N__17501;
    wire N__17494;
    wire N__17493;
    wire N__17492;
    wire N__17485;
    wire N__17484;
    wire N__17483;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17450;
    wire N__17449;
    wire N__17448;
    wire N__17447;
    wire N__17444;
    wire N__17443;
    wire N__17442;
    wire N__17439;
    wire N__17436;
    wire N__17431;
    wire N__17428;
    wire N__17423;
    wire N__17422;
    wire N__17421;
    wire N__17420;
    wire N__17419;
    wire N__17418;
    wire N__17417;
    wire N__17416;
    wire N__17415;
    wire N__17412;
    wire N__17409;
    wire N__17406;
    wire N__17401;
    wire N__17400;
    wire N__17397;
    wire N__17394;
    wire N__17393;
    wire N__17390;
    wire N__17379;
    wire N__17370;
    wire N__17363;
    wire N__17360;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17342;
    wire N__17339;
    wire N__17336;
    wire N__17335;
    wire N__17332;
    wire N__17331;
    wire N__17330;
    wire N__17329;
    wire N__17328;
    wire N__17327;
    wire N__17326;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17318;
    wire N__17317;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17303;
    wire N__17300;
    wire N__17299;
    wire N__17294;
    wire N__17289;
    wire N__17284;
    wire N__17281;
    wire N__17272;
    wire N__17269;
    wire N__17256;
    wire N__17255;
    wire N__17254;
    wire N__17253;
    wire N__17252;
    wire N__17249;
    wire N__17248;
    wire N__17247;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17239;
    wire N__17238;
    wire N__17237;
    wire N__17234;
    wire N__17225;
    wire N__17220;
    wire N__17217;
    wire N__17214;
    wire N__17211;
    wire N__17210;
    wire N__17209;
    wire N__17206;
    wire N__17201;
    wire N__17198;
    wire N__17193;
    wire N__17186;
    wire N__17183;
    wire N__17178;
    wire N__17169;
    wire N__17166;
    wire N__17165;
    wire N__17164;
    wire N__17159;
    wire N__17156;
    wire N__17151;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17115;
    wire N__17114;
    wire N__17113;
    wire N__17112;
    wire N__17111;
    wire N__17110;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17094;
    wire N__17093;
    wire N__17086;
    wire N__17081;
    wire N__17080;
    wire N__17079;
    wire N__17074;
    wire N__17069;
    wire N__17064;
    wire N__17063;
    wire N__17062;
    wire N__17061;
    wire N__17058;
    wire N__17055;
    wire N__17054;
    wire N__17051;
    wire N__17050;
    wire N__17049;
    wire N__17046;
    wire N__17045;
    wire N__17044;
    wire N__17043;
    wire N__17040;
    wire N__17035;
    wire N__17032;
    wire N__17027;
    wire N__17024;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17006;
    wire N__17005;
    wire N__17004;
    wire N__17003;
    wire N__17002;
    wire N__16991;
    wire N__16982;
    wire N__16977;
    wire N__16974;
    wire N__16971;
    wire N__16970;
    wire N__16967;
    wire N__16966;
    wire N__16965;
    wire N__16964;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16939;
    wire N__16938;
    wire N__16933;
    wire N__16932;
    wire N__16931;
    wire N__16930;
    wire N__16929;
    wire N__16928;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16893;
    wire N__16890;
    wire N__16875;
    wire N__16874;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16866;
    wire N__16865;
    wire N__16864;
    wire N__16863;
    wire N__16862;
    wire N__16861;
    wire N__16860;
    wire N__16859;
    wire N__16856;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16848;
    wire N__16845;
    wire N__16842;
    wire N__16841;
    wire N__16840;
    wire N__16837;
    wire N__16826;
    wire N__16821;
    wire N__16816;
    wire N__16813;
    wire N__16802;
    wire N__16799;
    wire N__16788;
    wire N__16785;
    wire N__16784;
    wire N__16783;
    wire N__16782;
    wire N__16781;
    wire N__16780;
    wire N__16777;
    wire N__16774;
    wire N__16771;
    wire N__16768;
    wire N__16767;
    wire N__16764;
    wire N__16761;
    wire N__16758;
    wire N__16755;
    wire N__16754;
    wire N__16751;
    wire N__16744;
    wire N__16743;
    wire N__16742;
    wire N__16741;
    wire N__16738;
    wire N__16733;
    wire N__16730;
    wire N__16725;
    wire N__16722;
    wire N__16721;
    wire N__16720;
    wire N__16717;
    wire N__16716;
    wire N__16713;
    wire N__16708;
    wire N__16703;
    wire N__16692;
    wire N__16683;
    wire N__16682;
    wire N__16681;
    wire N__16678;
    wire N__16675;
    wire N__16674;
    wire N__16673;
    wire N__16672;
    wire N__16671;
    wire N__16670;
    wire N__16669;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16661;
    wire N__16660;
    wire N__16659;
    wire N__16658;
    wire N__16657;
    wire N__16656;
    wire N__16653;
    wire N__16642;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16630;
    wire N__16627;
    wire N__16616;
    wire N__16611;
    wire N__16596;
    wire N__16595;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16570;
    wire N__16569;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16553;
    wire N__16548;
    wire N__16547;
    wire N__16546;
    wire N__16543;
    wire N__16542;
    wire N__16541;
    wire N__16538;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16512;
    wire N__16509;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16473;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16465;
    wire N__16464;
    wire N__16463;
    wire N__16460;
    wire N__16459;
    wire N__16458;
    wire N__16455;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16433;
    wire N__16422;
    wire N__16421;
    wire N__16418;
    wire N__16417;
    wire N__16416;
    wire N__16415;
    wire N__16414;
    wire N__16413;
    wire N__16410;
    wire N__16409;
    wire N__16406;
    wire N__16403;
    wire N__16398;
    wire N__16393;
    wire N__16390;
    wire N__16387;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16365;
    wire N__16364;
    wire N__16363;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16347;
    wire N__16346;
    wire N__16345;
    wire N__16344;
    wire N__16343;
    wire N__16342;
    wire N__16337;
    wire N__16334;
    wire N__16329;
    wire N__16320;
    wire N__16311;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16289;
    wire N__16288;
    wire N__16287;
    wire N__16286;
    wire N__16285;
    wire N__16284;
    wire N__16283;
    wire N__16280;
    wire N__16279;
    wire N__16278;
    wire N__16269;
    wire N__16262;
    wire N__16259;
    wire N__16254;
    wire N__16253;
    wire N__16252;
    wire N__16251;
    wire N__16248;
    wire N__16245;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16218;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16202;
    wire N__16201;
    wire N__16200;
    wire N__16199;
    wire N__16194;
    wire N__16193;
    wire N__16188;
    wire N__16185;
    wire N__16184;
    wire N__16183;
    wire N__16180;
    wire N__16177;
    wire N__16176;
    wire N__16175;
    wire N__16172;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16153;
    wire N__16152;
    wire N__16147;
    wire N__16144;
    wire N__16137;
    wire N__16136;
    wire N__16135;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16115;
    wire N__16104;
    wire N__16103;
    wire N__16102;
    wire N__16099;
    wire N__16098;
    wire N__16097;
    wire N__16096;
    wire N__16095;
    wire N__16094;
    wire N__16093;
    wire N__16092;
    wire N__16091;
    wire N__16090;
    wire N__16087;
    wire N__16084;
    wire N__16083;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16066;
    wire N__16065;
    wire N__16060;
    wire N__16059;
    wire N__16058;
    wire N__16057;
    wire N__16056;
    wire N__16055;
    wire N__16054;
    wire N__16053;
    wire N__16050;
    wire N__16049;
    wire N__16046;
    wire N__16045;
    wire N__16042;
    wire N__16037;
    wire N__16032;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16014;
    wire N__16011;
    wire N__16006;
    wire N__16001;
    wire N__15994;
    wire N__15989;
    wire N__15984;
    wire N__15981;
    wire N__15978;
    wire N__15971;
    wire N__15964;
    wire N__15945;
    wire N__15944;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15928;
    wire N__15921;
    wire N__15920;
    wire N__15919;
    wire N__15918;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15906;
    wire N__15903;
    wire N__15902;
    wire N__15901;
    wire N__15900;
    wire N__15899;
    wire N__15898;
    wire N__15897;
    wire N__15896;
    wire N__15895;
    wire N__15894;
    wire N__15893;
    wire N__15892;
    wire N__15891;
    wire N__15890;
    wire N__15889;
    wire N__15888;
    wire N__15887;
    wire N__15886;
    wire N__15885;
    wire N__15884;
    wire N__15883;
    wire N__15882;
    wire N__15881;
    wire N__15880;
    wire N__15879;
    wire N__15878;
    wire N__15877;
    wire N__15876;
    wire N__15875;
    wire N__15874;
    wire N__15873;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15863;
    wire N__15860;
    wire N__15859;
    wire N__15858;
    wire N__15857;
    wire N__15856;
    wire N__15855;
    wire N__15854;
    wire N__15853;
    wire N__15852;
    wire N__15851;
    wire N__15850;
    wire N__15849;
    wire N__15848;
    wire N__15753;
    wire N__15750;
    wire N__15747;
    wire N__15744;
    wire N__15741;
    wire N__15738;
    wire N__15735;
    wire N__15734;
    wire N__15733;
    wire N__15732;
    wire N__15731;
    wire N__15730;
    wire N__15729;
    wire N__15726;
    wire N__15725;
    wire N__15716;
    wire N__15715;
    wire N__15714;
    wire N__15713;
    wire N__15708;
    wire N__15705;
    wire N__15702;
    wire N__15699;
    wire N__15692;
    wire N__15691;
    wire N__15690;
    wire N__15689;
    wire N__15686;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15668;
    wire N__15665;
    wire N__15654;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15646;
    wire N__15643;
    wire N__15642;
    wire N__15641;
    wire N__15640;
    wire N__15639;
    wire N__15638;
    wire N__15637;
    wire N__15636;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15628;
    wire N__15627;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15611;
    wire N__15610;
    wire N__15603;
    wire N__15598;
    wire N__15591;
    wire N__15584;
    wire N__15581;
    wire N__15570;
    wire N__15567;
    wire N__15564;
    wire N__15561;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15551;
    wire N__15548;
    wire N__15547;
    wire N__15546;
    wire N__15545;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15533;
    wire N__15532;
    wire N__15531;
    wire N__15530;
    wire N__15527;
    wire N__15526;
    wire N__15523;
    wire N__15520;
    wire N__15515;
    wire N__15510;
    wire N__15503;
    wire N__15492;
    wire N__15491;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15459;
    wire N__15458;
    wire N__15457;
    wire N__15456;
    wire N__15453;
    wire N__15452;
    wire N__15451;
    wire N__15450;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15442;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15432;
    wire N__15427;
    wire N__15426;
    wire N__15425;
    wire N__15422;
    wire N__15421;
    wire N__15420;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15398;
    wire N__15393;
    wire N__15386;
    wire N__15369;
    wire N__15368;
    wire N__15367;
    wire N__15366;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15347;
    wire N__15346;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15334;
    wire N__15331;
    wire N__15326;
    wire N__15321;
    wire N__15318;
    wire N__15309;
    wire N__15308;
    wire N__15307;
    wire N__15306;
    wire N__15305;
    wire N__15302;
    wire N__15301;
    wire N__15296;
    wire N__15293;
    wire N__15292;
    wire N__15291;
    wire N__15288;
    wire N__15283;
    wire N__15280;
    wire N__15275;
    wire N__15272;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15256;
    wire N__15249;
    wire N__15248;
    wire N__15247;
    wire N__15244;
    wire N__15241;
    wire N__15240;
    wire N__15237;
    wire N__15236;
    wire N__15235;
    wire N__15232;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15198;
    wire N__15195;
    wire N__15192;
    wire N__15189;
    wire N__15188;
    wire N__15187;
    wire N__15184;
    wire N__15183;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15168;
    wire N__15167;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15149;
    wire N__15138;
    wire N__15137;
    wire N__15136;
    wire N__15135;
    wire N__15134;
    wire N__15133;
    wire N__15132;
    wire N__15131;
    wire N__15130;
    wire N__15127;
    wire N__15120;
    wire N__15109;
    wire N__15102;
    wire N__15101;
    wire N__15100;
    wire N__15099;
    wire N__15096;
    wire N__15095;
    wire N__15092;
    wire N__15089;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15074;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15053;
    wire N__15052;
    wire N__15051;
    wire N__15050;
    wire N__15049;
    wire N__15048;
    wire N__15047;
    wire N__15046;
    wire N__15043;
    wire N__15034;
    wire N__15027;
    wire N__15018;
    wire N__15009;
    wire N__15006;
    wire N__15003;
    wire N__15002;
    wire N__15001;
    wire N__15000;
    wire N__14999;
    wire N__14998;
    wire N__14995;
    wire N__14994;
    wire N__14993;
    wire N__14992;
    wire N__14989;
    wire N__14988;
    wire N__14987;
    wire N__14984;
    wire N__14979;
    wire N__14976;
    wire N__14975;
    wire N__14972;
    wire N__14965;
    wire N__14962;
    wire N__14961;
    wire N__14958;
    wire N__14955;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14937;
    wire N__14934;
    wire N__14931;
    wire N__14928;
    wire N__14925;
    wire N__14918;
    wire N__14907;
    wire N__14906;
    wire N__14903;
    wire N__14902;
    wire N__14897;
    wire N__14896;
    wire N__14893;
    wire N__14892;
    wire N__14891;
    wire N__14890;
    wire N__14889;
    wire N__14888;
    wire N__14887;
    wire N__14884;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14870;
    wire N__14867;
    wire N__14866;
    wire N__14861;
    wire N__14856;
    wire N__14851;
    wire N__14848;
    wire N__14843;
    wire N__14832;
    wire N__14831;
    wire N__14828;
    wire N__14827;
    wire N__14826;
    wire N__14823;
    wire N__14822;
    wire N__14821;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14809;
    wire N__14806;
    wire N__14801;
    wire N__14796;
    wire N__14793;
    wire N__14792;
    wire N__14791;
    wire N__14790;
    wire N__14787;
    wire N__14780;
    wire N__14773;
    wire N__14766;
    wire N__14763;
    wire N__14760;
    wire N__14757;
    wire N__14754;
    wire N__14751;
    wire N__14750;
    wire N__14749;
    wire N__14748;
    wire N__14747;
    wire N__14746;
    wire N__14745;
    wire N__14744;
    wire N__14743;
    wire N__14738;
    wire N__14735;
    wire N__14734;
    wire N__14721;
    wire N__14720;
    wire N__14719;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14686;
    wire N__14679;
    wire N__14676;
    wire N__14675;
    wire N__14674;
    wire N__14673;
    wire N__14672;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14664;
    wire N__14661;
    wire N__14658;
    wire N__14655;
    wire N__14652;
    wire N__14651;
    wire N__14650;
    wire N__14647;
    wire N__14638;
    wire N__14637;
    wire N__14634;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14619;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14605;
    wire N__14602;
    wire N__14597;
    wire N__14592;
    wire N__14587;
    wire N__14580;
    wire N__14577;
    wire N__14574;
    wire N__14573;
    wire N__14572;
    wire N__14569;
    wire N__14568;
    wire N__14565;
    wire N__14562;
    wire N__14559;
    wire N__14558;
    wire N__14557;
    wire N__14556;
    wire N__14555;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14537;
    wire N__14530;
    wire N__14527;
    wire N__14514;
    wire N__14511;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14503;
    wire N__14502;
    wire N__14501;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14484;
    wire N__14481;
    wire N__14472;
    wire N__14469;
    wire N__14466;
    wire N__14463;
    wire N__14462;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14454;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14439;
    wire N__14434;
    wire N__14427;
    wire N__14426;
    wire N__14425;
    wire N__14422;
    wire N__14417;
    wire N__14416;
    wire N__14415;
    wire N__14410;
    wire N__14405;
    wire N__14400;
    wire N__14399;
    wire N__14398;
    wire N__14397;
    wire N__14392;
    wire N__14387;
    wire N__14386;
    wire N__14385;
    wire N__14384;
    wire N__14381;
    wire N__14378;
    wire N__14373;
    wire N__14370;
    wire N__14369;
    wire N__14366;
    wire N__14363;
    wire N__14360;
    wire N__14355;
    wire N__14346;
    wire N__14343;
    wire N__14340;
    wire N__14337;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14322;
    wire N__14319;
    wire N__14316;
    wire N__14313;
    wire N__14312;
    wire N__14309;
    wire N__14308;
    wire N__14307;
    wire N__14306;
    wire N__14303;
    wire N__14300;
    wire N__14295;
    wire N__14292;
    wire N__14289;
    wire N__14288;
    wire N__14287;
    wire N__14286;
    wire N__14285;
    wire N__14284;
    wire N__14279;
    wire N__14274;
    wire N__14271;
    wire N__14262;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14235;
    wire N__14234;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14223;
    wire N__14222;
    wire N__14221;
    wire N__14214;
    wire N__14209;
    wire N__14206;
    wire N__14199;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14191;
    wire N__14190;
    wire N__14189;
    wire N__14188;
    wire N__14187;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14171;
    wire N__14168;
    wire N__14167;
    wire N__14162;
    wire N__14161;
    wire N__14160;
    wire N__14159;
    wire N__14158;
    wire N__14155;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14135;
    wire N__14130;
    wire N__14121;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14113;
    wire N__14112;
    wire N__14111;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14091;
    wire N__14090;
    wire N__14089;
    wire N__14088;
    wire N__14083;
    wire N__14080;
    wire N__14075;
    wire N__14072;
    wire N__14071;
    wire N__14070;
    wire N__14067;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14048;
    wire N__14043;
    wire N__14036;
    wire N__14033;
    wire N__14028;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__14012;
    wire N__14011;
    wire N__14010;
    wire N__14007;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13997;
    wire N__13996;
    wire N__13995;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13973;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13929;
    wire N__13926;
    wire N__13925;
    wire N__13920;
    wire N__13919;
    wire N__13918;
    wire N__13917;
    wire N__13916;
    wire N__13915;
    wire N__13914;
    wire N__13913;
    wire N__13910;
    wire N__13903;
    wire N__13900;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13866;
    wire N__13857;
    wire N__13856;
    wire N__13853;
    wire N__13852;
    wire N__13851;
    wire N__13848;
    wire N__13847;
    wire N__13844;
    wire N__13843;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13828;
    wire N__13827;
    wire N__13826;
    wire N__13823;
    wire N__13822;
    wire N__13813;
    wire N__13808;
    wire N__13805;
    wire N__13800;
    wire N__13791;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13781;
    wire N__13780;
    wire N__13779;
    wire N__13776;
    wire N__13775;
    wire N__13772;
    wire N__13771;
    wire N__13770;
    wire N__13769;
    wire N__13766;
    wire N__13765;
    wire N__13764;
    wire N__13763;
    wire N__13762;
    wire N__13759;
    wire N__13758;
    wire N__13757;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13737;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13718;
    wire N__13715;
    wire N__13708;
    wire N__13705;
    wire N__13694;
    wire N__13683;
    wire N__13680;
    wire N__13679;
    wire N__13676;
    wire N__13673;
    wire N__13668;
    wire N__13665;
    wire N__13662;
    wire N__13659;
    wire N__13656;
    wire N__13655;
    wire N__13654;
    wire N__13649;
    wire N__13646;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13615;
    wire N__13612;
    wire N__13609;
    wire N__13606;
    wire N__13599;
    wire N__13596;
    wire N__13593;
    wire N__13592;
    wire N__13589;
    wire N__13586;
    wire N__13581;
    wire N__13578;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13570;
    wire N__13567;
    wire N__13564;
    wire N__13561;
    wire N__13554;
    wire N__13551;
    wire N__13548;
    wire N__13547;
    wire N__13546;
    wire N__13545;
    wire N__13544;
    wire N__13543;
    wire N__13542;
    wire N__13541;
    wire N__13540;
    wire N__13539;
    wire N__13538;
    wire N__13537;
    wire N__13536;
    wire N__13535;
    wire N__13534;
    wire N__13533;
    wire N__13532;
    wire N__13531;
    wire N__13530;
    wire N__13529;
    wire N__13528;
    wire N__13527;
    wire N__13526;
    wire N__13525;
    wire N__13524;
    wire N__13523;
    wire N__13522;
    wire N__13521;
    wire N__13520;
    wire N__13519;
    wire N__13518;
    wire N__13517;
    wire N__13516;
    wire N__13515;
    wire N__13514;
    wire N__13513;
    wire N__13512;
    wire N__13511;
    wire N__13510;
    wire N__13509;
    wire N__13508;
    wire N__13507;
    wire N__13506;
    wire N__13505;
    wire N__13504;
    wire N__13503;
    wire N__13502;
    wire N__13501;
    wire N__13500;
    wire N__13499;
    wire N__13498;
    wire N__13497;
    wire N__13496;
    wire N__13495;
    wire N__13494;
    wire N__13493;
    wire N__13492;
    wire N__13491;
    wire N__13490;
    wire N__13489;
    wire N__13488;
    wire N__13487;
    wire N__13486;
    wire N__13485;
    wire N__13484;
    wire N__13483;
    wire N__13350;
    wire N__13347;
    wire N__13344;
    wire N__13341;
    wire N__13338;
    wire N__13335;
    wire N__13334;
    wire N__13331;
    wire N__13328;
    wire N__13323;
    wire N__13322;
    wire N__13321;
    wire N__13318;
    wire N__13313;
    wire N__13308;
    wire N__13307;
    wire N__13306;
    wire N__13303;
    wire N__13298;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13278;
    wire N__13275;
    wire N__13272;
    wire N__13269;
    wire N__13266;
    wire N__13263;
    wire N__13260;
    wire N__13257;
    wire N__13254;
    wire N__13251;
    wire N__13248;
    wire N__13245;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13233;
    wire N__13230;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13218;
    wire N__13215;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13184;
    wire N__13183;
    wire N__13180;
    wire N__13179;
    wire N__13178;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13161;
    wire N__13152;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13133;
    wire N__13130;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13116;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13086;
    wire N__13083;
    wire N__13082;
    wire N__13081;
    wire N__13078;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13070;
    wire N__13069;
    wire N__13066;
    wire N__13061;
    wire N__13060;
    wire N__13057;
    wire N__13052;
    wire N__13047;
    wire N__13044;
    wire N__13035;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__12999;
    wire N__12996;
    wire N__12993;
    wire N__12990;
    wire N__12989;
    wire N__12988;
    wire N__12987;
    wire N__12986;
    wire N__12985;
    wire N__12980;
    wire N__12977;
    wire N__12970;
    wire N__12963;
    wire N__12962;
    wire N__12961;
    wire N__12958;
    wire N__12955;
    wire N__12954;
    wire N__12953;
    wire N__12952;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12935;
    wire N__12924;
    wire N__12921;
    wire N__12918;
    wire N__12917;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12872;
    wire N__12869;
    wire N__12868;
    wire N__12865;
    wire N__12862;
    wire N__12859;
    wire N__12856;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12839;
    wire N__12838;
    wire N__12837;
    wire N__12836;
    wire N__12835;
    wire N__12834;
    wire N__12831;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12819;
    wire N__12814;
    wire N__12813;
    wire N__12812;
    wire N__12811;
    wire N__12810;
    wire N__12805;
    wire N__12800;
    wire N__12799;
    wire N__12798;
    wire N__12797;
    wire N__12796;
    wire N__12795;
    wire N__12794;
    wire N__12791;
    wire N__12788;
    wire N__12779;
    wire N__12774;
    wire N__12767;
    wire N__12764;
    wire N__12761;
    wire N__12758;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12731;
    wire N__12730;
    wire N__12729;
    wire N__12728;
    wire N__12727;
    wire N__12724;
    wire N__12719;
    wire N__12716;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12704;
    wire N__12699;
    wire N__12694;
    wire N__12691;
    wire N__12686;
    wire N__12681;
    wire N__12678;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12651;
    wire N__12648;
    wire N__12645;
    wire N__12644;
    wire N__12643;
    wire N__12640;
    wire N__12635;
    wire N__12632;
    wire N__12631;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12619;
    wire N__12618;
    wire N__12617;
    wire N__12614;
    wire N__12609;
    wire N__12604;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12582;
    wire N__12579;
    wire N__12576;
    wire N__12575;
    wire N__12572;
    wire N__12571;
    wire N__12570;
    wire N__12569;
    wire N__12566;
    wire N__12565;
    wire N__12564;
    wire N__12563;
    wire N__12562;
    wire N__12561;
    wire N__12558;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12540;
    wire N__12535;
    wire N__12534;
    wire N__12531;
    wire N__12528;
    wire N__12525;
    wire N__12524;
    wire N__12523;
    wire N__12516;
    wire N__12513;
    wire N__12510;
    wire N__12505;
    wire N__12500;
    wire N__12497;
    wire N__12486;
    wire N__12483;
    wire N__12482;
    wire N__12479;
    wire N__12478;
    wire N__12477;
    wire N__12476;
    wire N__12475;
    wire N__12472;
    wire N__12471;
    wire N__12470;
    wire N__12469;
    wire N__12468;
    wire N__12467;
    wire N__12466;
    wire N__12463;
    wire N__12462;
    wire N__12461;
    wire N__12460;
    wire N__12451;
    wire N__12448;
    wire N__12445;
    wire N__12440;
    wire N__12433;
    wire N__12430;
    wire N__12429;
    wire N__12428;
    wire N__12427;
    wire N__12426;
    wire N__12425;
    wire N__12424;
    wire N__12421;
    wire N__12420;
    wire N__12415;
    wire N__12412;
    wire N__12405;
    wire N__12400;
    wire N__12399;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12379;
    wire N__12376;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12360;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12338;
    wire N__12337;
    wire N__12334;
    wire N__12329;
    wire N__12324;
    wire N__12323;
    wire N__12322;
    wire N__12317;
    wire N__12316;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12294;
    wire N__12293;
    wire N__12292;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12276;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12252;
    wire N__12249;
    wire N__12246;
    wire N__12243;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12231;
    wire N__12230;
    wire N__12229;
    wire N__12226;
    wire N__12225;
    wire N__12224;
    wire N__12223;
    wire N__12222;
    wire N__12217;
    wire N__12214;
    wire N__12213;
    wire N__12212;
    wire N__12209;
    wire N__12204;
    wire N__12201;
    wire N__12198;
    wire N__12195;
    wire N__12192;
    wire N__12187;
    wire N__12182;
    wire N__12181;
    wire N__12178;
    wire N__12173;
    wire N__12168;
    wire N__12165;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12131;
    wire N__12130;
    wire N__12127;
    wire N__12124;
    wire N__12119;
    wire N__12114;
    wire N__12113;
    wire N__12112;
    wire N__12105;
    wire N__12102;
    wire N__12101;
    wire N__12098;
    wire N__12097;
    wire N__12094;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12078;
    wire N__12077;
    wire N__12076;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12064;
    wire N__12061;
    wire N__12054;
    wire N__12053;
    wire N__12052;
    wire N__12049;
    wire N__12048;
    wire N__12041;
    wire N__12040;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12028;
    wire N__12021;
    wire N__12018;
    wire N__12017;
    wire N__12016;
    wire N__12013;
    wire N__12010;
    wire N__12009;
    wire N__12008;
    wire N__12007;
    wire N__12006;
    wire N__12003;
    wire N__11998;
    wire N__11995;
    wire N__11986;
    wire N__11979;
    wire N__11978;
    wire N__11977;
    wire N__11976;
    wire N__11975;
    wire N__11972;
    wire N__11967;
    wire N__11962;
    wire N__11955;
    wire N__11954;
    wire N__11953;
    wire N__11952;
    wire N__11949;
    wire N__11946;
    wire N__11943;
    wire N__11940;
    wire N__11937;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11921;
    wire N__11920;
    wire N__11919;
    wire N__11918;
    wire N__11915;
    wire N__11914;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11893;
    wire N__11880;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11849;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11841;
    wire N__11836;
    wire N__11831;
    wire N__11826;
    wire N__11825;
    wire N__11824;
    wire N__11823;
    wire N__11822;
    wire N__11821;
    wire N__11812;
    wire N__11807;
    wire N__11802;
    wire N__11799;
    wire N__11798;
    wire N__11797;
    wire N__11792;
    wire N__11789;
    wire N__11784;
    wire N__11783;
    wire N__11782;
    wire N__11781;
    wire N__11780;
    wire N__11771;
    wire N__11768;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11699;
    wire N__11698;
    wire N__11695;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11687;
    wire N__11686;
    wire N__11685;
    wire N__11684;
    wire N__11683;
    wire N__11680;
    wire N__11677;
    wire N__11674;
    wire N__11671;
    wire N__11664;
    wire N__11663;
    wire N__11662;
    wire N__11661;
    wire N__11658;
    wire N__11655;
    wire N__11652;
    wire N__11649;
    wire N__11642;
    wire N__11631;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11613;
    wire N__11610;
    wire N__11607;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11599;
    wire N__11598;
    wire N__11597;
    wire N__11596;
    wire N__11595;
    wire N__11590;
    wire N__11589;
    wire N__11588;
    wire N__11587;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11562;
    wire N__11557;
    wire N__11544;
    wire N__11541;
    wire N__11538;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11520;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11478;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11435;
    wire N__11432;
    wire N__11429;
    wire N__11426;
    wire N__11423;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11341;
    wire N__11336;
    wire N__11333;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11319;
    wire N__11316;
    wire N__11315;
    wire N__11314;
    wire N__11311;
    wire N__11306;
    wire N__11305;
    wire N__11304;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11283;
    wire N__11280;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11256;
    wire N__11255;
    wire N__11254;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11242;
    wire N__11235;
    wire N__11234;
    wire N__11233;
    wire N__11232;
    wire N__11229;
    wire N__11228;
    wire N__11227;
    wire N__11226;
    wire N__11225;
    wire N__11224;
    wire N__11223;
    wire N__11222;
    wire N__11221;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11193;
    wire N__11192;
    wire N__11191;
    wire N__11190;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11177;
    wire N__11170;
    wire N__11167;
    wire N__11166;
    wire N__11165;
    wire N__11164;
    wire N__11163;
    wire N__11162;
    wire N__11159;
    wire N__11150;
    wire N__11147;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11120;
    wire N__11109;
    wire N__11106;
    wire N__11105;
    wire N__11104;
    wire N__11103;
    wire N__11100;
    wire N__11095;
    wire N__11092;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11076;
    wire N__11073;
    wire N__11072;
    wire N__11071;
    wire N__11070;
    wire N__11069;
    wire N__11068;
    wire N__11065;
    wire N__11058;
    wire N__11053;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11045;
    wire N__11044;
    wire N__11043;
    wire N__11042;
    wire N__11041;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11025;
    wire N__11018;
    wire N__11013;
    wire N__11008;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10959;
    wire N__10956;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10941;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10920;
    wire N__10917;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10907;
    wire N__10906;
    wire N__10905;
    wire N__10896;
    wire N__10893;
    wire N__10892;
    wire N__10891;
    wire N__10884;
    wire N__10881;
    wire N__10880;
    wire N__10879;
    wire N__10878;
    wire N__10877;
    wire N__10876;
    wire N__10873;
    wire N__10868;
    wire N__10861;
    wire N__10854;
    wire N__10851;
    wire N__10850;
    wire N__10849;
    wire N__10848;
    wire N__10839;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10824;
    wire N__10823;
    wire N__10818;
    wire N__10815;
    wire N__10814;
    wire N__10813;
    wire N__10812;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10790;
    wire N__10785;
    wire N__10776;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10761;
    wire N__10758;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10748;
    wire N__10745;
    wire N__10744;
    wire N__10741;
    wire N__10736;
    wire N__10731;
    wire N__10730;
    wire N__10727;
    wire N__10726;
    wire N__10719;
    wire N__10716;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10701;
    wire N__10700;
    wire N__10697;
    wire N__10696;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10684;
    wire N__10677;
    wire N__10674;
    wire N__10673;
    wire N__10672;
    wire N__10671;
    wire N__10670;
    wire N__10669;
    wire N__10668;
    wire N__10667;
    wire N__10666;
    wire N__10663;
    wire N__10656;
    wire N__10651;
    wire N__10644;
    wire N__10641;
    wire N__10632;
    wire N__10629;
    wire N__10626;
    wire N__10623;
    wire N__10620;
    wire N__10617;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10584;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10548;
    wire N__10547;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10532;
    wire N__10527;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10506;
    wire N__10503;
    wire N__10500;
    wire N__10497;
    wire N__10494;
    wire N__10491;
    wire N__10488;
    wire N__10485;
    wire N__10482;
    wire N__10479;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10434;
    wire N__10431;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10418;
    wire N__10415;
    wire N__10414;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10400;
    wire N__10395;
    wire N__10392;
    wire N__10389;
    wire N__10386;
    wire N__10383;
    wire N__10380;
    wire N__10377;
    wire N__10374;
    wire N__10371;
    wire N__10370;
    wire N__10369;
    wire N__10366;
    wire N__10365;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10350;
    wire N__10347;
    wire N__10344;
    wire N__10339;
    wire N__10336;
    wire N__10333;
    wire N__10330;
    wire N__10325;
    wire N__10320;
    wire N__10317;
    wire N__10316;
    wire N__10313;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10298;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10266;
    wire N__10263;
    wire N__10262;
    wire N__10257;
    wire N__10254;
    wire N__10251;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10226;
    wire N__10225;
    wire N__10224;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10197;
    wire N__10196;
    wire N__10195;
    wire N__10192;
    wire N__10187;
    wire N__10184;
    wire N__10183;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10171;
    wire N__10164;
    wire N__10163;
    wire N__10160;
    wire N__10159;
    wire N__10156;
    wire N__10155;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10135;
    wire N__10128;
    wire N__10127;
    wire N__10124;
    wire N__10119;
    wire N__10116;
    wire N__10115;
    wire N__10114;
    wire N__10113;
    wire N__10112;
    wire N__10111;
    wire N__10106;
    wire N__10105;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10074;
    wire N__10073;
    wire N__10072;
    wire N__10071;
    wire N__10070;
    wire N__10069;
    wire N__10064;
    wire N__10063;
    wire N__10060;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10032;
    wire N__10031;
    wire N__10030;
    wire N__10027;
    wire N__10024;
    wire N__10023;
    wire N__10020;
    wire N__10015;
    wire N__10014;
    wire N__10013;
    wire N__10010;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9991;
    wire N__9988;
    wire N__9985;
    wire N__9972;
    wire N__9971;
    wire N__9970;
    wire N__9969;
    wire N__9964;
    wire N__9961;
    wire N__9958;
    wire N__9955;
    wire N__9952;
    wire N__9945;
    wire N__9944;
    wire N__9939;
    wire N__9936;
    wire N__9935;
    wire N__9934;
    wire N__9931;
    wire N__9930;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9912;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9900;
    wire N__9897;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9889;
    wire N__9888;
    wire N__9885;
    wire N__9880;
    wire N__9879;
    wire N__9876;
    wire N__9875;
    wire N__9874;
    wire N__9873;
    wire N__9872;
    wire N__9871;
    wire N__9870;
    wire N__9865;
    wire N__9862;
    wire N__9853;
    wire N__9846;
    wire N__9845;
    wire N__9842;
    wire N__9835;
    wire N__9832;
    wire N__9825;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9791;
    wire N__9790;
    wire N__9785;
    wire N__9782;
    wire N__9777;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9765;
    wire N__9762;
    wire N__9761;
    wire N__9760;
    wire N__9759;
    wire N__9756;
    wire N__9749;
    wire N__9746;
    wire N__9741;
    wire N__9738;
    wire N__9735;
    wire N__9732;
    wire N__9731;
    wire N__9730;
    wire N__9727;
    wire N__9722;
    wire N__9717;
    wire N__9714;
    wire N__9713;
    wire N__9710;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9690;
    wire N__9687;
    wire N__9686;
    wire N__9683;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9671;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9659;
    wire N__9658;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9635;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9618;
    wire N__9615;
    wire N__9614;
    wire N__9611;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9591;
    wire N__9588;
    wire N__9585;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9573;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9540;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9528;
    wire N__9527;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9515;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9497;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9485;
    wire N__9480;
    wire N__9477;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9462;
    wire N__9459;
    wire N__9458;
    wire N__9453;
    wire N__9450;
    wire N__9449;
    wire N__9446;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9431;
    wire N__9430;
    wire N__9429;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9411;
    wire N__9410;
    wire N__9407;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9390;
    wire N__9387;
    wire N__9384;
    wire N__9381;
    wire N__9378;
    wire N__9375;
    wire N__9372;
    wire N__9371;
    wire N__9370;
    wire N__9367;
    wire N__9366;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9351;
    wire N__9342;
    wire N__9339;
    wire N__9336;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9323;
    wire N__9322;
    wire N__9319;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9304;
    wire N__9297;
    wire N__9294;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9282;
    wire N__9279;
    wire N__9276;
    wire N__9273;
    wire N__9270;
    wire N__9267;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9236;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9228;
    wire N__9221;
    wire N__9218;
    wire N__9217;
    wire N__9212;
    wire N__9209;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9138;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9083;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9048;
    wire N__9047;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9036;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9021;
    wire N__9018;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8990;
    wire N__8989;
    wire N__8988;
    wire N__8987;
    wire N__8984;
    wire N__8979;
    wire N__8974;
    wire N__8971;
    wire N__8964;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8927;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8919;
    wire N__8918;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8886;
    wire N__8885;
    wire N__8882;
    wire N__8881;
    wire N__8880;
    wire N__8879;
    wire N__8876;
    wire N__8867;
    wire N__8862;
    wire N__8859;
    wire N__8858;
    wire N__8857;
    wire N__8854;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8842;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8820;
    wire N__8817;
    wire N__8816;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8808;
    wire N__8805;
    wire N__8800;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8774;
    wire N__8773;
    wire N__8772;
    wire N__8769;
    wire N__8766;
    wire N__8761;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8745;
    wire N__8744;
    wire N__8743;
    wire N__8742;
    wire N__8741;
    wire N__8738;
    wire N__8737;
    wire N__8732;
    wire N__8731;
    wire N__8730;
    wire N__8729;
    wire N__8728;
    wire N__8727;
    wire N__8726;
    wire N__8725;
    wire N__8724;
    wire N__8723;
    wire N__8722;
    wire N__8721;
    wire N__8718;
    wire N__8715;
    wire N__8710;
    wire N__8707;
    wire N__8700;
    wire N__8693;
    wire N__8682;
    wire N__8667;
    wire N__8666;
    wire N__8665;
    wire N__8664;
    wire N__8661;
    wire N__8660;
    wire N__8659;
    wire N__8658;
    wire N__8657;
    wire N__8656;
    wire N__8655;
    wire N__8654;
    wire N__8653;
    wire N__8652;
    wire N__8651;
    wire N__8650;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8628;
    wire N__8625;
    wire N__8620;
    wire N__8613;
    wire N__8606;
    wire N__8599;
    wire N__8580;
    wire N__8577;
    wire N__8576;
    wire N__8575;
    wire N__8574;
    wire N__8571;
    wire N__8570;
    wire N__8569;
    wire N__8568;
    wire N__8567;
    wire N__8566;
    wire N__8565;
    wire N__8564;
    wire N__8563;
    wire N__8562;
    wire N__8561;
    wire N__8560;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8536;
    wire N__8529;
    wire N__8522;
    wire N__8519;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8492;
    wire N__8491;
    wire N__8488;
    wire N__8483;
    wire N__8478;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8454;
    wire N__8451;
    wire N__8450;
    wire N__8445;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8426;
    wire N__8425;
    wire N__8422;
    wire N__8417;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8405;
    wire N__8404;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8392;
    wire N__8385;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8334;
    wire N__8331;
    wire N__8328;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8316;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8256;
    wire N__8253;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8141;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8129;
    wire N__8124;
    wire N__8121;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8100;
    wire N__8097;
    wire N__8096;
    wire N__8095;
    wire N__8094;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8083;
    wire N__8082;
    wire N__8077;
    wire N__8074;
    wire N__8065;
    wire N__8058;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8028;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7962;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7940;
    wire N__7939;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7927;
    wire N__7920;
    wire N__7919;
    wire N__7918;
    wire N__7915;
    wire N__7914;
    wire N__7911;
    wire N__7908;
    wire N__7905;
    wire N__7904;
    wire N__7899;
    wire N__7894;
    wire N__7891;
    wire N__7884;
    wire N__7881;
    wire N__7878;
    wire N__7875;
    wire N__7872;
    wire N__7871;
    wire N__7870;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7858;
    wire N__7851;
    wire N__7848;
    wire N__7847;
    wire N__7846;
    wire N__7845;
    wire N__7840;
    wire N__7835;
    wire N__7830;
    wire N__7827;
    wire N__7824;
    wire N__7823;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7813;
    wire N__7806;
    wire N__7803;
    wire N__7802;
    wire N__7801;
    wire N__7798;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7784;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7733;
    wire N__7730;
    wire N__7727;
    wire N__7726;
    wire N__7721;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7704;
    wire N__7703;
    wire N__7702;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7690;
    wire N__7683;
    wire N__7682;
    wire N__7677;
    wire N__7676;
    wire N__7675;
    wire N__7674;
    wire N__7673;
    wire N__7672;
    wire N__7671;
    wire N__7670;
    wire N__7667;
    wire N__7662;
    wire N__7659;
    wire N__7654;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7646;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7587;
    wire N__7586;
    wire N__7585;
    wire N__7584;
    wire N__7583;
    wire N__7582;
    wire N__7581;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7556;
    wire N__7555;
    wire N__7554;
    wire N__7553;
    wire N__7546;
    wire N__7541;
    wire N__7540;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7517;
    wire N__7516;
    wire N__7515;
    wire N__7512;
    wire N__7507;
    wire N__7504;
    wire N__7497;
    wire N__7494;
    wire N__7493;
    wire N__7490;
    wire N__7489;
    wire N__7488;
    wire N__7485;
    wire N__7484;
    wire N__7483;
    wire N__7480;
    wire N__7477;
    wire N__7474;
    wire N__7471;
    wire N__7466;
    wire N__7457;
    wire N__7452;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7444;
    wire N__7441;
    wire N__7440;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7425;
    wire N__7422;
    wire N__7413;
    wire N__7412;
    wire N__7411;
    wire N__7408;
    wire N__7403;
    wire N__7400;
    wire N__7395;
    wire N__7394;
    wire N__7391;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7378;
    wire N__7371;
    wire N__7368;
    wire N__7367;
    wire N__7364;
    wire N__7363;
    wire N__7360;
    wire N__7357;
    wire N__7354;
    wire N__7347;
    wire N__7344;
    wire N__7343;
    wire N__7342;
    wire N__7341;
    wire N__7338;
    wire N__7335;
    wire N__7330;
    wire N__7327;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7310;
    wire N__7307;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7295;
    wire N__7290;
    wire N__7289;
    wire N__7288;
    wire N__7285;
    wire N__7282;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7263;
    wire N__7262;
    wire N__7259;
    wire N__7258;
    wire N__7257;
    wire N__7254;
    wire N__7251;
    wire N__7246;
    wire N__7243;
    wire N__7240;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7196;
    wire N__7195;
    wire N__7194;
    wire N__7193;
    wire N__7192;
    wire N__7191;
    wire N__7190;
    wire N__7189;
    wire N__7180;
    wire N__7169;
    wire N__7164;
    wire N__7161;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7143;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7133;
    wire N__7132;
    wire N__7131;
    wire N__7130;
    wire N__7129;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7101;
    wire N__7100;
    wire N__7099;
    wire N__7096;
    wire N__7095;
    wire N__7094;
    wire N__7089;
    wire N__7086;
    wire N__7083;
    wire N__7080;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7052;
    wire N__7049;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7019;
    wire N__7016;
    wire N__7015;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7003;
    wire N__6996;
    wire N__6993;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6968;
    wire N__6967;
    wire N__6966;
    wire N__6963;
    wire N__6958;
    wire N__6955;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6941;
    wire N__6936;
    wire N__6933;
    wire N__6932;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6879;
    wire N__6878;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6815;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6801;
    wire N__6798;
    wire N__6797;
    wire N__6796;
    wire N__6793;
    wire N__6792;
    wire N__6785;
    wire N__6782;
    wire N__6777;
    wire N__6776;
    wire N__6775;
    wire N__6774;
    wire N__6773;
    wire N__6762;
    wire N__6759;
    wire N__6758;
    wire N__6757;
    wire N__6756;
    wire N__6753;
    wire N__6748;
    wire N__6745;
    wire N__6738;
    wire N__6737;
    wire N__6736;
    wire N__6735;
    wire N__6732;
    wire N__6723;
    wire N__6720;
    wire N__6719;
    wire N__6718;
    wire N__6717;
    wire N__6716;
    wire N__6707;
    wire N__6704;
    wire N__6699;
    wire N__6696;
    wire N__6695;
    wire N__6694;
    wire N__6691;
    wire N__6686;
    wire N__6685;
    wire N__6680;
    wire N__6677;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6644;
    wire N__6643;
    wire N__6642;
    wire N__6639;
    wire N__6636;
    wire N__6633;
    wire N__6632;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6609;
    wire N__6606;
    wire N__6605;
    wire N__6604;
    wire N__6603;
    wire N__6600;
    wire N__6593;
    wire N__6588;
    wire N__6587;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6573;
    wire N__6570;
    wire N__6569;
    wire N__6568;
    wire N__6565;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6553;
    wire N__6546;
    wire N__6545;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6479;
    wire N__6478;
    wire N__6477;
    wire N__6476;
    wire N__6473;
    wire N__6464;
    wire N__6459;
    wire N__6458;
    wire N__6457;
    wire N__6456;
    wire N__6455;
    wire N__6452;
    wire N__6447;
    wire N__6442;
    wire N__6435;
    wire N__6432;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6420;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6366;
    wire N__6363;
    wire N__6362;
    wire N__6359;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6336;
    wire N__6333;
    wire N__6330;
    wire clk_in_c;
    wire GNDG0;
    wire VCCG0;
    wire \Lab_UT.secuu0.un131_ci_3_cascade_ ;
    wire \Lab_UT.secuu0.un142_ci_0 ;
    wire \Lab_UT.secuu0.un131_ci_3 ;
    wire \Lab_UT.secuu0.un87_ci ;
    wire \Lab_UT.secuu0.un87_ci_cascade_ ;
    wire Lab_UT_L3_tx_data_0_4_cascade_;
    wire Lab_UT_dspStr_un29_dOut_0_cascade_;
    wire bfn_1_8_0_;
    wire \Lab_UT.dspStr.un1_cnt_3_cry_0 ;
    wire \Lab_UT.dspStr.un1_cnt_3_cry_1 ;
    wire \Lab_UT.dspStr.un1_cnt_3_cry_2 ;
    wire \uu2.un1_w_user_lfZ0Z_4 ;
    wire L3_tx_data_0_cascade_;
    wire \uu2.un1_w_user_lf_0 ;
    wire \uu2.un1_w_user_lf_0_cascade_ ;
    wire \INVuu2.w_addr_user_4C_net ;
    wire uart_RXD;
    wire \uu2.un447_ci_3_cascade_ ;
    wire \uu2.o_adder_vbuf_w_addr_user_7 ;
    wire \uu2.mem0.w_addr_6 ;
    wire \uu2.mem0.w_addr_7 ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire \uu2.un447_ci_3 ;
    wire \uu2.vbuf_w_addr_user.un469_ci_0_cascade_ ;
    wire \uu2.o_adder_vbuf_w_addr_user_8 ;
    wire \Lab_UT.secuu0.un230_ci_1 ;
    wire \Lab_UT.secuu0.un109_ci ;
    wire \Lab_UT.secuu0.un197_ci_9_cascade_ ;
    wire \Lab_UT.secuu0.l_countZ0Z_14 ;
    wire \Lab_UT.secuu0.l_countZ0Z_15 ;
    wire \Lab_UT.secuu0.l_countZ0Z_4 ;
    wire \Lab_UT.secuu0.l_countZ0Z_5 ;
    wire \Lab_UT.secuu0.l_precountZ0Z_3 ;
    wire \Lab_UT.secuu0.l_countZ0Z_1 ;
    wire \Lab_UT.secuu0.l_precountZ0Z_1 ;
    wire \Lab_UT.secuu0.l_countZ0Z_2 ;
    wire \Lab_UT.secuu0.l_precountZ0Z_2 ;
    wire \Lab_UT.secuu0.l_countZ0Z_0 ;
    wire \Lab_UT.secuu0.un4_l_count_14_cascade_ ;
    wire \Lab_UT.secuu0.un4_l_count_0_8 ;
    wire \Lab_UT.secuu0.un4_l_count_12 ;
    wire \Lab_UT.secuu0.un4_l_count_13 ;
    wire \Lab_UT.secuu0.un4_l_count_18_cascade_ ;
    wire \Lab_UT.dspStr.cnt11_1_cascade_ ;
    wire \Lab_UT.dspStr.cnt11_0_i ;
    wire \Lab_UT.secuu0.un11_l_count_i ;
    wire Lab_UT_dspStr_un29_dOut_0;
    wire \uu2.un27_w_addr_user_0 ;
    wire \Lab_UT.dspStr.cntZ0Z_0 ;
    wire \uu2.un1_w_user_lfZ0Z_1 ;
    wire \uu2.un1_w_user_lfZ0Z_3 ;
    wire \uu2.un1_w_user_cr_0_0 ;
    wire \uu2.un1_w_user_crZ0Z_2 ;
    wire L3_tx_data_rdy;
    wire \uu2.un1_w_user_crZ0Z_2_cascade_ ;
    wire \uu2.un19_w_addr_userZ0Z_0_cascade_ ;
    wire L3_tx_data_7;
    wire \uu2.mem0.w_data_7 ;
    wire \uu2.un1_w_user_cr_5Z0Z_1 ;
    wire Lab_UT_L3_tx_data_2_0_cascade_;
    wire \uu2.un1_w_user_crZ0Z_5 ;
    wire Lab_UT_L3_tx_data_0_6;
    wire \uu2.mem0.w_data_6 ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \uu2.mem0.w_addr_8 ;
    wire Lab_UT_L3_tx_data_2_0;
    wire \uu2.mem0.w_addr_1 ;
    wire L3_tx_data_2;
    wire \uu2.mem0.w_data_2 ;
    wire \uu2.un2_w_addr_user_5_cascade_ ;
    wire \uu2.un2_w_addr_user_4 ;
    wire \uu2.un2_w_addr_user ;
    wire \uu2.un27_w_addr_user_i ;
    wire \INVuu2.w_addr_user_3C_net ;
    wire \uu2.w_addr_user_RNIKHHELZ0Z_2 ;
    wire \uu2.o_adder_vbuf_w_addr_user_3 ;
    wire \uu2.w_addr_userZ0Z_1 ;
    wire \uu2.un425_ci ;
    wire \uu2.r_data_wire_3 ;
    wire \Lab_UT.secuu0.l_countZ0Z_10 ;
    wire \Lab_UT.secuu0.un186_ci_0_cascade_ ;
    wire \Lab_UT.secuu0.l_countZ0Z_8 ;
    wire \Lab_UT.secuu0.l_countZ0Z_9 ;
    wire \Lab_UT.secuu0.l_countZ0Z_7 ;
    wire \Lab_UT.secuu0.l_countZ0Z_3 ;
    wire \Lab_UT.secuu0.l_countZ0Z_11 ;
    wire \Lab_UT.secuu0.un4_l_count_11_cascade_ ;
    wire \Lab_UT.secuu0.l_countZ0Z_6 ;
    wire \Lab_UT.secuu0.un4_l_count_16 ;
    wire \Lab_UT.secuu0.l_countZ0Z_17 ;
    wire \Lab_UT.secuu0.un241_ci_2 ;
    wire \Lab_UT.secuu0.l_countZ0Z_16 ;
    wire \Lab_UT.secuu0.un263_ci ;
    wire \Lab_UT.secuu0.l_countZ0Z_18 ;
    wire \Lab_UT.secuu0.un197_ci_9 ;
    wire \Lab_UT.secuu0.l_countZ0Z_12 ;
    wire \Lab_UT.secuu0.un153_ci ;
    wire \Lab_UT.secuu0.un208_ci_0 ;
    wire \Lab_UT.secuu0.l_countZ0Z_13 ;
    wire \Lab_UT.secuu0.un11_l_count_i_g ;
    wire \Lab_UT.secuu0.l_precountZ0Z_0 ;
    wire \uu2.un425_ci_0_cascade_ ;
    wire \uu2.vbuf_raddr.un469_ci_0_cascade_ ;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.r_addrZ0Z_5 ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \uu2.vbuf_raddr.un447_ci_3 ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.vbuf_raddr.un447_ci_3_cascade_ ;
    wire \uu2.un425_ci_0 ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_21 ;
    wire \uu2.mem0.w_data_0 ;
    wire \uu2.mem0.w_data_ns_1_5 ;
    wire \uu2.mem0.w_data_5 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_17 ;
    wire \uu2.mem0.G_14_0_a6_0_cascade_ ;
    wire \uu2.mem0.N_7_0_cascade_ ;
    wire \uu2.mem0.w_data_1 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_22 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_ ;
    wire \uu2.mem0.w_data_4 ;
    wire \uu2.mem0.G_14_0_a6_0_0_1 ;
    wire \uu2.mem0.w_data_3 ;
    wire \uu2.N_326_0_cascade_ ;
    wire \uu2.bitmap_pmux_1_1_a8_1_2_0 ;
    wire \uu2.N_326_0 ;
    wire \uu2.bitmap_pmux_1_1_a8_1_1_cascade_ ;
    wire \uu2.bitmap_pmux_1_1_a8_0_1 ;
    wire \uu2.bitmap_pmux_1_1_1_tz ;
    wire \uu2.bitmap_pmux_1_1_1_tz_cascade_ ;
    wire L3_tx_data_3;
    wire \uu2.mem0.w_data_1_0_0_3 ;
    wire latticehx1k_pll_inst_PLLOUTCORE_i;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.mem0.w_addr_0 ;
    wire \INVuu2.w_addr_displaying_1C_net ;
    wire \uu2.r_data_wire_1 ;
    wire \uu2.r_data_wire_2 ;
    wire \uu2.r_data_wire_0 ;
    wire \uu2.r_data_wire_4 ;
    wire \uu2.r_data_wire_5 ;
    wire \uu2.r_data_wire_6 ;
    wire \uu2.r_data_wire_7 ;
    wire vbuf_tx_data_0;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire vbuf_tx_data_1;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire vbuf_tx_data_2;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire vbuf_tx_data_3;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire vbuf_tx_data_4;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire vbuf_tx_data_5;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire bfn_5_3_0_;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \buart.Z_rx.N_144_cascade_ ;
    wire buart__rx_bitcount_4;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire buart__rx_bitcount_1;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire CONSTANT_ONE_NET;
    wire \resetGen.reset_count_2_i_0_a3_5Z0Z_4_cascade_ ;
    wire bu_rx_data_5;
    wire \resetGen.reset_count_2_i_0_a3_6Z0Z_4 ;
    wire \resetGen.reset_count_2_i_0_a3_4Z0Z_4 ;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire \buart.Z_rx.N_129_cascade_ ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire \buart.Z_rx.N_39 ;
    wire Lab_UT_rx_data_4;
    wire Lab_UT_rx_data_3;
    wire \Lab_UT.dictrluu0.N_103_1_cascade_ ;
    wire Lab_UT_rx_data_5;
    wire \uu2.un1_w_user_lf_3Z0Z_1 ;
    wire Lab_UT_dspStr_cnt_1;
    wire Lab_UT_dspStr_cnt_3;
    wire \uu2.mem0.N_26_1_cascade_ ;
    wire Lab_UT_dspStr_cnt_2;
    wire \Lab_UT.Lab3U00.bu_rx_data_rdy_0 ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.mem0.w_addr_2 ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.mem0.w_addr_3 ;
    wire \uu2.mem0.G_14_0_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_32_cascade_ ;
    wire \uu2.mem0.G_14_0_1 ;
    wire \uu2.N_329_0_cascade_ ;
    wire \uu2.Z_decfrac105_7 ;
    wire N_52_0;
    wire L3_segment2_0_0;
    wire \uu2.mem0.N_2159_0_cascade_ ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_20 ;
    wire L3_segment2_0;
    wire \uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4_cascade_ ;
    wire \uu2.mem0.g2_0 ;
    wire \uu2.mem0.N_5_cascade_ ;
    wire \uu2.mem0.bitmap_pmux_1_1_0_0 ;
    wire \uu2.mem0.N_14 ;
    wire \uu2.mem0.N_18 ;
    wire \uu2.mem0.un1_segment3_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_34 ;
    wire \uu2.Z_decfrac106 ;
    wire \uu2.mem0.un1_segment3_m2_1 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_47_cascade_ ;
    wire \uu2.mem0.un1_segment3_1_1 ;
    wire \uu2.mem0.N_2160_0 ;
    wire N_52;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_48 ;
    wire vbuf_tx_data_6;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire vbuf_tx_data_7;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire \uu2.mem0.w_addr_4 ;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \uu2.mem0.w_addr_5 ;
    wire \uu2.Z_decfrac106_2 ;
    wire \uu2.mem0.N_2160_1 ;
    wire bfn_6_1_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire bfn_6_3_0_;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \buart.Z_rx.ser_clk_cascade_ ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire bu_rx_data_7;
    wire bu_rx_data_6;
    wire bu_rx_data_2;
    wire bu_rx_data_4;
    wire bu_rx_data_3;
    wire Lab_UT_rx_data_7;
    wire Lab_UT_rx_data_1;
    wire Lab_UT_rx_data_6;
    wire \Lab_UT.rx_data_rdy ;
    wire buart__rx_bitcount_0;
    wire buart__rx_bitcount_2;
    wire buart__rx_bitcount_3;
    wire N_118;
    wire bu_rx_data_rdy;
    wire \buart.Z_rx.ser_clk ;
    wire \buart.Z_rx.N_129 ;
    wire bu_rx_data_rdy_cascade_;
    wire \buart.Z_rx.startbit ;
    wire \buart.Z_rx.bitcount_e_0_RNII0231Z0Z_0 ;
    wire Lab_UT_dec3_segmentUQ_0_6_cascade_;
    wire N_71;
    wire N_71_cascade_;
    wire Lab_UT_dec3_segmentUQ_1_1_cascade_;
    wire \uu2.Z_decfrac105_7_2 ;
    wire \Lab_UT.rx_data_0 ;
    wire \Lab_UT.rx_dataZ0Z_2 ;
    wire \Lab_UT.dictrluu0.N_103_1 ;
    wire \Lab_UT.dicSelectLEDdisp ;
    wire \Lab_UT.dicSelectLEDdisp_cascade_ ;
    wire \Lab_UT.dictrluu0.N_72 ;
    wire \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_o2_2 ;
    wire \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_3 ;
    wire \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_4 ;
    wire \Lab_UT.dictrluu0.dicfsm.N_102_cascade_ ;
    wire \uu2.N_93 ;
    wire \uu2.N_49_cascade_ ;
    wire \uu2.un1_segment3_m4_s_2 ;
    wire \uu2.g0_i_o4_0_1 ;
    wire \uu2.un1_segment3_m4_ns_1 ;
    wire \uu2.g0_i_o4_3_cascade_ ;
    wire \uu2.un1_segment3_m4 ;
    wire \uu2.w_addr_displaying_4_rep1_RNIMMRIAZ0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_53_cascade_ ;
    wire \uu2.mem0.un1_segment3_1_2 ;
    wire \uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4 ;
    wire \uu2.mem0.un1_segment3_m2_2 ;
    wire \uu2.mem0.un1_segment3_m2_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_42_cascade_ ;
    wire \uu2.mem0.un1_segment3_1_0 ;
    wire \Lab_UT.didpuu0.didpmtens.q_5_0_0_2 ;
    wire \uu2.un1_segment4_1_amZ0 ;
    wire \uu2.un1_segment4_1_bmZ0_cascade_ ;
    wire \uu2.w_addr_displaying_fast_RNIPN54Z0Z_8_cascade_ ;
    wire \uu2.N_292 ;
    wire \uu2.un1_segment4_5_amZ0Z_1 ;
    wire \uu2.w_addr_displaying_fast_RNIV5694Z0Z_2 ;
    wire \uu2.N_290_0_i_0_cascade_ ;
    wire \uu2.w_addr_displaying_RNI362A1Z0Z_3 ;
    wire \uu2.un1_w_addr_displaying_19_cascade_ ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_ ;
    wire \uu2.mem0.N_5_0 ;
    wire \uu2.un1_segment3_s_0 ;
    wire \INVuu2.w_addr_displaying_5C_net ;
    wire \uu2.un1_segment4_5_bmZ0 ;
    wire \Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMUZ0Z_0_cascade_ ;
    wire led_c_2;
    wire \Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJZ0Z_0 ;
    wire bfn_7_2_0_;
    wire \buart.Z_tx.un1_bitcount_cry_0 ;
    wire \buart.Z_tx.un1_bitcount_cry_1 ;
    wire \buart.Z_tx.un1_bitcount_axb_3 ;
    wire \buart.Z_tx.un1_bitcount_cry_2 ;
    wire \buart.Z_tx.bitcount_RNIM5O32Z0Z_2 ;
    wire \buart.Z_tx.bitcount_RNIL4O32Z0Z_1 ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire buart__tx_uart_busy_0_cascade_;
    wire \buart.Z_tx.ser_clk ;
    wire \buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0 ;
    wire \resetGen.N_117 ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire \resetGen.N_117_cascade_ ;
    wire rst;
    wire \resetGen.reset_countZ0Z_0 ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \resetGen.reset_countZ0Z_4 ;
    wire \resetGen.N_96_cascade_ ;
    wire \resetGen.N_133 ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire buart__tx_uart_busy_0;
    wire vbuf_tx_data_rdy_cascade_;
    wire \uu2.vbuf_tx_data_rdy_0 ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \uu2.r_addrZ0Z_0 ;
    wire vbuf_tx_data_rdy;
    wire \uu2.r_addrZ0Z_2 ;
    wire \Lab_UT.secuu0.un4_l_count_0 ;
    wire \Lab_UT.secuu0.delay_lineZ0Z_0 ;
    wire \Lab_UT.secuu0.delay_lineZ0Z_1 ;
    wire \Lab_UT.didpuu0.didpmtens.N_122 ;
    wire N_84_cascade_;
    wire N_7;
    wire \uu2.un1_segment4_0_bmZ0 ;
    wire \uu2.un1_segment4_0_amZ0_cascade_ ;
    wire \uu2.un1_segment4_2_bmZ0 ;
    wire \uu2.un1_segment4_8_ns_1_cascade_ ;
    wire \uu2.un1_segment4_2_amZ0 ;
    wire \uu2.N_286 ;
    wire \Lab_UT.N_10_cascade_ ;
    wire \uu2.g0_i_o4_0_a8_2_2_cascade_ ;
    wire \uu2.w_addr_displaying_5_rep1_RNIVO2EZ0Z1 ;
    wire \uu2.N_315_1_0 ;
    wire \INVuu2.w_addr_displaying_fast_4C_net ;
    wire \uu2.N_94 ;
    wire \uu2.bitmap_pmux_1_1_3_tz_1_cascade_ ;
    wire \uu2.bitmap_pmux_1_1_3_tz ;
    wire \uu2.N_111_cascade_ ;
    wire \INVuu2.w_addr_displaying_4C_net ;
    wire \uu2.un1_segment4_sn_N_36_mux_0_cascade_ ;
    wire \uu2.gZ0Z1 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_54 ;
    wire \uu2.un1_segment4_sn_N_58_0 ;
    wire \uu2.N_2150_0 ;
    wire \uu2.un1_segment4_sn_N_38_0_0 ;
    wire \uu2.g2_1_cascade_ ;
    wire \uu2.N_299_0 ;
    wire \uu2.un1_w_addr_displaying_inv_4_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_43 ;
    wire \uu2.segment3_m_1Z0Z_6_cascade_ ;
    wire \uu2.segment3_m_2_6_cascade_ ;
    wire \uu2.un1_segment4_4_bmZ0 ;
    wire \uu2.un1_segment4_4_amZ0_cascade_ ;
    wire \uu2.mem0.G_14_0_a6_2_1 ;
    wire \uu2.mem0.bitmap_pmux_1_1_2_tz_0 ;
    wire \uu2.bitmap_pmux_1_1_2_tz_1_0 ;
    wire \uu2.bitmap_pmux_1_1_2_tz_1_0_cascade_ ;
    wire \uu2.mem0.bitmap_pmux_1_1_2_tz_cascade_ ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_33 ;
    wire \INVuu2.w_addr_displaying_2C_net ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \uu2.w_addr_displaying_RNI8NHB1Z0Z_2_cascade_ ;
    wire \uu2.w_addr_displaying_RNI18582Z0Z_8 ;
    wire \uu2.l_countZ0Z_2 ;
    wire \uu2.l_countZ0Z_0 ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.un3_r_clk_en_7 ;
    wire \uu2.un3_r_clk_en_0_0_cascade_ ;
    wire \uu2.un3_r_clk_en_6 ;
    wire uu2_un3_r_clk_en_0_cascade_;
    wire \uu2.un349_ci_0 ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.vbuf_count.un382_ci_8_1 ;
    wire \uu2.l_countZ0Z_8 ;
    wire \uu2.l_countZ0Z_4 ;
    wire \uu2.un316_ci ;
    wire \uu2.l_countZ0Z_5 ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu2.un382_ci ;
    wire uu2_un3_r_clk_en_0;
    wire \uu2.l_countZ0Z_10 ;
    wire \Lab_UT.didpuu0.countEnMones_cascade_ ;
    wire \Lab_UT.didpuu0.didpmones.countEnMones_0 ;
    wire \Lab_UT.didpuu0.countEnStens_cascade_ ;
    wire \uu2.un1_segment4_2_amZ0Z_1 ;
    wire \uu2.w_addr_displaying_4_0_i_6_cascade_ ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \uu2.g0_i_o4_0_a8_3_1 ;
    wire \uu2.w_addr_displaying_4_0_i_fast_6 ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \uu2.un15_w_data_displaying_cascade_ ;
    wire \uu2.un19_w_addr_userZ0Z_0 ;
    wire \uu2.un21_w_addr_displaying_i_cascade_ ;
    wire \INVuu2.w_addr_displaying_6C_net ;
    wire \uu2.un15_w_data_displaying ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.w_addr_displaying_4_0_i_rep1_6 ;
    wire \uu2.w_addr_displaying_5_rep1_RNI3HMTZ0_cascade_ ;
    wire \INVuu2.w_addr_displaying_6_rep1C_net ;
    wire \uu2.un1_segment4_sn_N_61 ;
    wire \uu2.w_addr_displaying_fast_RNI6N2KZ0Z_5_cascade_ ;
    wire \uu2.w_addr_displaying_fast_RNID5QHZ0Z_5 ;
    wire \uu2.un1_segment4_sn_N_39_0 ;
    wire \uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4 ;
    wire \uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4_cascade_ ;
    wire \uu2.w_addr_displaying_RNILB202Z0Z_4 ;
    wire \uu2.N_92 ;
    wire \INVuu2.w_addr_displaying_fast_3C_net ;
    wire \uu2.w_addr_displaying_fast_RNIN0TSZ0Z_4 ;
    wire \uu2.w_addr_displaying_fastZ0Z_4 ;
    wire \uu2.w_addr_displaying_fastZ0Z_2 ;
    wire \uu2.N_10_0 ;
    wire \Lab_UT.didpuu0.didpsones.N_38 ;
    wire \Lab_UT.didpuu0.didpsones.N_32 ;
    wire Lab_UT_dec0_un137_segmentUQ;
    wire \uu2.segment1_m_2Z0Z_0_cascade_ ;
    wire \uu2.segment1_m_0_cascade_ ;
    wire \uu2.w_addr_displayingZ0Z_3 ;
    wire \uu2.segment3_m_6 ;
    wire \uu2.un1_segment1_iv_0_cascade_ ;
    wire \uu2.un1_segment1_0 ;
    wire \Lab_UT.didpuu0.didpstens.countEnStens_0 ;
    wire \uu2.un1_segment4_3_bmZ0 ;
    wire \uu2.un1_segment4_3_amZ0_cascade_ ;
    wire \uu2.un1_segment4_9_ns_1 ;
    wire \uu2.N_289_cascade_ ;
    wire \uu2.w_addr_displaying_fast_RNIFU9M8Z0Z_8 ;
    wire \uu2.w_addr_displaying_fastZ0Z_3 ;
    wire \uu2.N_1 ;
    wire \uu2.w_addr_displaying_4_rep1_RNIAVDBZ0Z_0 ;
    wire \uu2.w_addr_displaying_fast_RNIKFIEZ0Z_6 ;
    wire \Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMUZ0Z_0_cascade_ ;
    wire led_c_3;
    wire \Lab_UT.didpuu0.ledDisp00.selLed_RNI67CIZ0Z_0 ;
    wire \Lab_UT.un11_segmentUQ_1 ;
    wire \Lab_UT.didpuu0.countEnMtens_0_a4_0_cascade_ ;
    wire \Lab_UT.didpuu0.countEnMtens_0_a4_1 ;
    wire \Lab_UT.didpuu0.countEnMtens_0_a4_1_cascade_ ;
    wire \Lab_UT.didpuu0.countEnStens ;
    wire \Lab_UT.didpuu0.countEnMtens ;
    wire \Lab_UT.un152_segmentUQ_1 ;
    wire \Lab_UT.didpuu0.countEnMones ;
    wire \uu2.un1_segment3_m5_bmZ0 ;
    wire bu_rx_data_1;
    wire bu_rx_data_0;
    wire \buart.Z_rx.N_41_i ;
    wire clk_g;
    wire \Lab_UT.sec_clkD ;
    wire \Lab_UT.didpuu0.clkSecStrbZ0 ;
    wire L3_segment3_2;
    wire L3_segment2_4_cascade_;
    wire \uu2.segment2_m_1Z0Z_6 ;
    wire Lab_UT_di_Stens_2;
    wire Lab_UT_di_Stens_3;
    wire \uu2.un1_segment3_m5_amZ0 ;
    wire \uu2.N_290_0_i_0 ;
    wire \uu2.un436_ci ;
    wire \INVuu2.w_addr_displaying_4_rep1C_net ;
    wire \uu2.w_addr_displaying_8_repZ0Z1 ;
    wire \uu2.un1_w_addr_displaying_35_0 ;
    wire \uu2.w_addr_displayingZ0Z_4 ;
    wire \uu2.un1_w_addr_displaying_35_0_cascade_ ;
    wire \uu2.un1_w_addr_displaying_inv_2 ;
    wire \uu2.N_813_0_cascade_ ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_58 ;
    wire \uu2.w_addr_displaying_7_repZ0Z1 ;
    wire \uu2.w_addr_displaying_4_repZ0Z1 ;
    wire \uu2.un1_segment3_m4_s_2_1 ;
    wire Lab_UT_di_Sones_2;
    wire Lab_UT_di_Sones_3;
    wire \uu2.un1_segment3_m0 ;
    wire \uu2.w_addr_displaying_fastZ0Z_6 ;
    wire L3_segment1_3_cascade_;
    wire \uu2.w_addr_displaying_fastZ0Z_5 ;
    wire \uu2.w_addr_displaying_fast_RNIQD7R4Z0Z_5 ;
    wire \uu2.N_315_1 ;
    wire \uu2.w_addr_displaying_4_rep2_RNI75VMZ0 ;
    wire \uu2.un1_segment3_m5 ;
    wire \uu2.N_813_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_59 ;
    wire \uu2.segment2_m_2Z0Z_5 ;
    wire \uu2.segment2_m_5 ;
    wire \uu2.w_addr_displaying_0_repZ0Z1 ;
    wire \uu2.w_addr_displaying_fastZ0Z_7 ;
    wire \uu2.w_addr_displaying_4_rep2_RNI4S6JZ0 ;
    wire \uu2.w_addr_displaying_fast_RNIEDBMZ0Z_7_cascade_ ;
    wire \uu2.un1_segment4_sn_N_38_0 ;
    wire \uu2.w_addr_displaying_4_repZ0Z2 ;
    wire \uu2.N_111 ;
    wire \uu2.w_addr_displaying_3_repZ0Z1 ;
    wire \uu2.Z_decfrac106_6 ;
    wire \uu2.un15_w_data_displaying_5 ;
    wire \uu2.w_addr_displaying_fastZ0Z_8 ;
    wire \INVuu2.w_addr_displaying_0_rep1C_net ;
    wire L3_segment4_2_cascade_;
    wire \uu2.N_280 ;
    wire Lab_UT_di_Mtens_2;
    wire Lab_UT_di_Mtens_3;
    wire L3_segment4_4;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \INVuu2.w_addr_displaying_2_rep1C_net ;
    wire \uu2.un1_w_addr_displaying_46_1 ;
    wire \uu2.un1_w_addr_displaying_46_1_cascade_ ;
    wire \uu2.w_addr_displaying_RNI8U3D2Z0Z_0 ;
    wire \uu2.w_addr_displaying_5_repZ0Z1 ;
    wire \uu2.w_addr_displaying_6_repZ0Z1 ;
    wire \uu2.w_addr_displaying_2_repZ0Z1 ;
    wire \uu2.un1_w_addr_displaying_38_1 ;
    wire \uu2.segment3_m_3Z0Z_1 ;
    wire \uu2.un1_w_addr_displaying_38_1_cascade_ ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire \uu2.segment3_m_1 ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.un21_w_addr_displaying_i ;
    wire \uu2.w_addr_displaying_fastZ0Z_0 ;
    wire \INVuu2.w_addr_displaying_0C_net ;
    wire rst_g;
    wire \uu2.mem0.N_2160_2 ;
    wire Lab_UT_di_Sones_0;
    wire Lab_UT_di_Stens_0;
    wire \Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11Z0Z_0_cascade_ ;
    wire led_c_0;
    wire Lab_UT_di_Mtens_0;
    wire \Lab_UT.didpuu0.ledDisp00.selLed_RNINURJZ0Z_0 ;
    wire Lab_UT_di_Stens_1;
    wire Lab_UT_di_Sones_1;
    wire \Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11Z0Z_0_cascade_ ;
    wire \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_1 ;
    wire led_c_1;
    wire \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_0 ;
    wire Lab_UT_di_Mtens_1;
    wire \Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJZ0Z_0 ;
    wire Lab_UT_di_Mones_2;
    wire Lab_UT_di_Mones_1;
    wire Lab_UT_di_Mones_3;
    wire Lab_UT_di_Mones_0;
    wire \uu2.N_2160_1_0_0 ;
    wire Lab_UT_dicRun;
    wire Lab_UT_l_oneSecPluse;
    wire led_c_4;
    wire _gnd_net_;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(latticehx1k_pll_inst_PLLOUTCORE_i),
            .REFERENCECLK(N__6339),
            .RESETB(N__8370),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__7968,N__7830,N__7878,N__7950,N__7920,N__7806,N__11109,N__11322,N__11283}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__6996,N__6495,N__6510,N__9297,N__9342,N__8964,N__9009,N__6981,N__8058}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,N__6870,dangling_wire_29,N__7026,dangling_wire_30,N__7752,dangling_wire_31,N__7995,dangling_wire_32,N__7980,dangling_wire_33,N__6948,dangling_wire_34,N__8013,dangling_wire_35,N__7770}),
            .RCLKE(N__11235),
            .RCLK(N__13508),
            .RE(N__11232),
            .WCLKE(N__8121),
            .WCLK(N__13509),
            .WE(N__8120));
    IO_PAD led_obuf_4_iopad (
            .OE(N__17566),
            .DIN(N__17565),
            .DOUT(N__17564),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__17566),
            .PADOUT(N__17565),
            .PADIN(N__17564),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16500),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_1_iopad (
            .OE(N__17557),
            .DIN(N__17556),
            .DOUT(N__17555),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__17557),
            .PADOUT(N__17556),
            .PADIN(N__17555),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17127),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__17548),
            .DIN(N__17547),
            .DOUT(N__17546),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__17548),
            .PADOUT(N__17547),
            .PADIN(N__17546),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8232),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__17539),
            .DIN(N__17538),
            .DOUT(N__17537),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__17539),
            .PADOUT(N__17538),
            .PADIN(N__17537),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_2_iopad (
            .OE(N__17530),
            .DIN(N__17529),
            .DOUT(N__17528),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__17530),
            .PADOUT(N__17529),
            .PADIN(N__17528),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10611),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_3_iopad (
            .OE(N__17521),
            .DIN(N__17520),
            .DOUT(N__17519),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__17521),
            .PADOUT(N__17520),
            .PADIN(N__17519),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13263),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_0_iopad (
            .OE(N__17512),
            .DIN(N__17511),
            .DOUT(N__17510),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__17512),
            .PADOUT(N__17511),
            .PADIN(N__17510),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17463),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__17503),
            .DIN(N__17502),
            .DOUT(N__17501),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__17503),
            .PADOUT(N__17502),
            .PADIN(N__17501),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__13514),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__17494),
            .DIN(N__17493),
            .DOUT(N__17492),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__17494),
            .PADOUT(N__17493),
            .PADIN(N__17492),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__17485),
            .DIN(N__17484),
            .DOUT(N__17483),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__17485),
            .PADOUT(N__17484),
            .PADIN(N__17483),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__4248 (
            .O(N__17466),
            .I(\Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11Z0Z_0_cascade_ ));
    IoInMux I__4247 (
            .O(N__17463),
            .I(N__17460));
    LocalMux I__4246 (
            .O(N__17460),
            .I(N__17457));
    Span12Mux_s3_h I__4245 (
            .O(N__17457),
            .I(N__17454));
    Odrv12 I__4244 (
            .O(N__17454),
            .I(led_c_0));
    InMux I__4243 (
            .O(N__17451),
            .I(N__17444));
    InMux I__4242 (
            .O(N__17450),
            .I(N__17439));
    InMux I__4241 (
            .O(N__17449),
            .I(N__17436));
    InMux I__4240 (
            .O(N__17448),
            .I(N__17431));
    InMux I__4239 (
            .O(N__17447),
            .I(N__17431));
    LocalMux I__4238 (
            .O(N__17444),
            .I(N__17428));
    InMux I__4237 (
            .O(N__17443),
            .I(N__17423));
    InMux I__4236 (
            .O(N__17442),
            .I(N__17423));
    LocalMux I__4235 (
            .O(N__17439),
            .I(N__17412));
    LocalMux I__4234 (
            .O(N__17436),
            .I(N__17409));
    LocalMux I__4233 (
            .O(N__17431),
            .I(N__17406));
    Span4Mux_v I__4232 (
            .O(N__17428),
            .I(N__17401));
    LocalMux I__4231 (
            .O(N__17423),
            .I(N__17401));
    CascadeMux I__4230 (
            .O(N__17422),
            .I(N__17397));
    CascadeMux I__4229 (
            .O(N__17421),
            .I(N__17394));
    InMux I__4228 (
            .O(N__17420),
            .I(N__17390));
    InMux I__4227 (
            .O(N__17419),
            .I(N__17379));
    InMux I__4226 (
            .O(N__17418),
            .I(N__17379));
    InMux I__4225 (
            .O(N__17417),
            .I(N__17379));
    InMux I__4224 (
            .O(N__17416),
            .I(N__17379));
    InMux I__4223 (
            .O(N__17415),
            .I(N__17379));
    Span4Mux_h I__4222 (
            .O(N__17412),
            .I(N__17370));
    Span4Mux_v I__4221 (
            .O(N__17409),
            .I(N__17370));
    Span4Mux_v I__4220 (
            .O(N__17406),
            .I(N__17370));
    Span4Mux_v I__4219 (
            .O(N__17401),
            .I(N__17370));
    InMux I__4218 (
            .O(N__17400),
            .I(N__17363));
    InMux I__4217 (
            .O(N__17397),
            .I(N__17363));
    InMux I__4216 (
            .O(N__17394),
            .I(N__17363));
    InMux I__4215 (
            .O(N__17393),
            .I(N__17360));
    LocalMux I__4214 (
            .O(N__17390),
            .I(Lab_UT_di_Mtens_0));
    LocalMux I__4213 (
            .O(N__17379),
            .I(Lab_UT_di_Mtens_0));
    Odrv4 I__4212 (
            .O(N__17370),
            .I(Lab_UT_di_Mtens_0));
    LocalMux I__4211 (
            .O(N__17363),
            .I(Lab_UT_di_Mtens_0));
    LocalMux I__4210 (
            .O(N__17360),
            .I(Lab_UT_di_Mtens_0));
    InMux I__4209 (
            .O(N__17349),
            .I(N__17346));
    LocalMux I__4208 (
            .O(N__17346),
            .I(\Lab_UT.didpuu0.ledDisp00.selLed_RNINURJZ0Z_0 ));
    InMux I__4207 (
            .O(N__17343),
            .I(N__17339));
    InMux I__4206 (
            .O(N__17342),
            .I(N__17336));
    LocalMux I__4205 (
            .O(N__17339),
            .I(N__17332));
    LocalMux I__4204 (
            .O(N__17336),
            .I(N__17322));
    InMux I__4203 (
            .O(N__17335),
            .I(N__17319));
    Span4Mux_h I__4202 (
            .O(N__17332),
            .I(N__17313));
    InMux I__4201 (
            .O(N__17331),
            .I(N__17310));
    InMux I__4200 (
            .O(N__17330),
            .I(N__17303));
    InMux I__4199 (
            .O(N__17329),
            .I(N__17303));
    InMux I__4198 (
            .O(N__17328),
            .I(N__17303));
    InMux I__4197 (
            .O(N__17327),
            .I(N__17300));
    InMux I__4196 (
            .O(N__17326),
            .I(N__17294));
    InMux I__4195 (
            .O(N__17325),
            .I(N__17294));
    Span4Mux_v I__4194 (
            .O(N__17322),
            .I(N__17289));
    LocalMux I__4193 (
            .O(N__17319),
            .I(N__17289));
    InMux I__4192 (
            .O(N__17318),
            .I(N__17284));
    InMux I__4191 (
            .O(N__17317),
            .I(N__17284));
    InMux I__4190 (
            .O(N__17316),
            .I(N__17281));
    Sp12to4 I__4189 (
            .O(N__17313),
            .I(N__17272));
    LocalMux I__4188 (
            .O(N__17310),
            .I(N__17272));
    LocalMux I__4187 (
            .O(N__17303),
            .I(N__17272));
    LocalMux I__4186 (
            .O(N__17300),
            .I(N__17272));
    InMux I__4185 (
            .O(N__17299),
            .I(N__17269));
    LocalMux I__4184 (
            .O(N__17294),
            .I(Lab_UT_di_Stens_1));
    Odrv4 I__4183 (
            .O(N__17289),
            .I(Lab_UT_di_Stens_1));
    LocalMux I__4182 (
            .O(N__17284),
            .I(Lab_UT_di_Stens_1));
    LocalMux I__4181 (
            .O(N__17281),
            .I(Lab_UT_di_Stens_1));
    Odrv12 I__4180 (
            .O(N__17272),
            .I(Lab_UT_di_Stens_1));
    LocalMux I__4179 (
            .O(N__17269),
            .I(Lab_UT_di_Stens_1));
    CascadeMux I__4178 (
            .O(N__17256),
            .I(N__17249));
    CascadeMux I__4177 (
            .O(N__17255),
            .I(N__17243));
    InMux I__4176 (
            .O(N__17254),
            .I(N__17240));
    InMux I__4175 (
            .O(N__17253),
            .I(N__17234));
    InMux I__4174 (
            .O(N__17252),
            .I(N__17225));
    InMux I__4173 (
            .O(N__17249),
            .I(N__17225));
    InMux I__4172 (
            .O(N__17248),
            .I(N__17225));
    InMux I__4171 (
            .O(N__17247),
            .I(N__17225));
    InMux I__4170 (
            .O(N__17246),
            .I(N__17220));
    InMux I__4169 (
            .O(N__17243),
            .I(N__17220));
    LocalMux I__4168 (
            .O(N__17240),
            .I(N__17217));
    InMux I__4167 (
            .O(N__17239),
            .I(N__17214));
    CascadeMux I__4166 (
            .O(N__17238),
            .I(N__17211));
    InMux I__4165 (
            .O(N__17237),
            .I(N__17206));
    LocalMux I__4164 (
            .O(N__17234),
            .I(N__17201));
    LocalMux I__4163 (
            .O(N__17225),
            .I(N__17201));
    LocalMux I__4162 (
            .O(N__17220),
            .I(N__17198));
    Span4Mux_v I__4161 (
            .O(N__17217),
            .I(N__17193));
    LocalMux I__4160 (
            .O(N__17214),
            .I(N__17193));
    InMux I__4159 (
            .O(N__17211),
            .I(N__17186));
    InMux I__4158 (
            .O(N__17210),
            .I(N__17186));
    InMux I__4157 (
            .O(N__17209),
            .I(N__17186));
    LocalMux I__4156 (
            .O(N__17206),
            .I(N__17183));
    Span4Mux_v I__4155 (
            .O(N__17201),
            .I(N__17178));
    Span4Mux_v I__4154 (
            .O(N__17198),
            .I(N__17178));
    Odrv4 I__4153 (
            .O(N__17193),
            .I(Lab_UT_di_Sones_1));
    LocalMux I__4152 (
            .O(N__17186),
            .I(Lab_UT_di_Sones_1));
    Odrv12 I__4151 (
            .O(N__17183),
            .I(Lab_UT_di_Sones_1));
    Odrv4 I__4150 (
            .O(N__17178),
            .I(Lab_UT_di_Sones_1));
    CascadeMux I__4149 (
            .O(N__17169),
            .I(\Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11Z0Z_0_cascade_ ));
    InMux I__4148 (
            .O(N__17166),
            .I(N__17159));
    InMux I__4147 (
            .O(N__17165),
            .I(N__17159));
    InMux I__4146 (
            .O(N__17164),
            .I(N__17156));
    LocalMux I__4145 (
            .O(N__17159),
            .I(N__17151));
    LocalMux I__4144 (
            .O(N__17156),
            .I(N__17151));
    Span4Mux_h I__4143 (
            .O(N__17151),
            .I(N__17147));
    InMux I__4142 (
            .O(N__17150),
            .I(N__17144));
    Span4Mux_v I__4141 (
            .O(N__17147),
            .I(N__17140));
    LocalMux I__4140 (
            .O(N__17144),
            .I(N__17137));
    InMux I__4139 (
            .O(N__17143),
            .I(N__17134));
    Odrv4 I__4138 (
            .O(N__17140),
            .I(\Lab_UT.didpuu0.ledDisp00.selLedZ0Z_1 ));
    Odrv12 I__4137 (
            .O(N__17137),
            .I(\Lab_UT.didpuu0.ledDisp00.selLedZ0Z_1 ));
    LocalMux I__4136 (
            .O(N__17134),
            .I(\Lab_UT.didpuu0.ledDisp00.selLedZ0Z_1 ));
    IoInMux I__4135 (
            .O(N__17127),
            .I(N__17124));
    LocalMux I__4134 (
            .O(N__17124),
            .I(N__17121));
    Span4Mux_s3_h I__4133 (
            .O(N__17121),
            .I(N__17118));
    Odrv4 I__4132 (
            .O(N__17118),
            .I(led_c_1));
    InMux I__4131 (
            .O(N__17115),
            .I(N__17101));
    InMux I__4130 (
            .O(N__17114),
            .I(N__17101));
    InMux I__4129 (
            .O(N__17113),
            .I(N__17101));
    InMux I__4128 (
            .O(N__17112),
            .I(N__17101));
    InMux I__4127 (
            .O(N__17111),
            .I(N__17098));
    InMux I__4126 (
            .O(N__17110),
            .I(N__17095));
    LocalMux I__4125 (
            .O(N__17101),
            .I(N__17086));
    LocalMux I__4124 (
            .O(N__17098),
            .I(N__17086));
    LocalMux I__4123 (
            .O(N__17095),
            .I(N__17086));
    InMux I__4122 (
            .O(N__17094),
            .I(N__17081));
    InMux I__4121 (
            .O(N__17093),
            .I(N__17081));
    Span12Mux_s6_h I__4120 (
            .O(N__17086),
            .I(N__17074));
    LocalMux I__4119 (
            .O(N__17081),
            .I(N__17074));
    InMux I__4118 (
            .O(N__17080),
            .I(N__17069));
    InMux I__4117 (
            .O(N__17079),
            .I(N__17069));
    Odrv12 I__4116 (
            .O(N__17074),
            .I(\Lab_UT.didpuu0.ledDisp00.selLedZ0Z_0 ));
    LocalMux I__4115 (
            .O(N__17069),
            .I(\Lab_UT.didpuu0.ledDisp00.selLedZ0Z_0 ));
    InMux I__4114 (
            .O(N__17064),
            .I(N__17058));
    CascadeMux I__4113 (
            .O(N__17063),
            .I(N__17055));
    InMux I__4112 (
            .O(N__17062),
            .I(N__17051));
    InMux I__4111 (
            .O(N__17061),
            .I(N__17046));
    LocalMux I__4110 (
            .O(N__17058),
            .I(N__17040));
    InMux I__4109 (
            .O(N__17055),
            .I(N__17035));
    InMux I__4108 (
            .O(N__17054),
            .I(N__17035));
    LocalMux I__4107 (
            .O(N__17051),
            .I(N__17032));
    InMux I__4106 (
            .O(N__17050),
            .I(N__17027));
    InMux I__4105 (
            .O(N__17049),
            .I(N__17027));
    LocalMux I__4104 (
            .O(N__17046),
            .I(N__17024));
    InMux I__4103 (
            .O(N__17045),
            .I(N__17017));
    InMux I__4102 (
            .O(N__17044),
            .I(N__17017));
    InMux I__4101 (
            .O(N__17043),
            .I(N__17017));
    Span4Mux_v I__4100 (
            .O(N__17040),
            .I(N__17014));
    LocalMux I__4099 (
            .O(N__17035),
            .I(N__17011));
    Span4Mux_v I__4098 (
            .O(N__17032),
            .I(N__17006));
    LocalMux I__4097 (
            .O(N__17027),
            .I(N__17006));
    Span4Mux_v I__4096 (
            .O(N__17024),
            .I(N__16991));
    LocalMux I__4095 (
            .O(N__17017),
            .I(N__16991));
    Span4Mux_h I__4094 (
            .O(N__17014),
            .I(N__16991));
    Span4Mux_v I__4093 (
            .O(N__17011),
            .I(N__16991));
    Span4Mux_v I__4092 (
            .O(N__17006),
            .I(N__16991));
    InMux I__4091 (
            .O(N__17005),
            .I(N__16982));
    InMux I__4090 (
            .O(N__17004),
            .I(N__16982));
    InMux I__4089 (
            .O(N__17003),
            .I(N__16982));
    InMux I__4088 (
            .O(N__17002),
            .I(N__16982));
    Odrv4 I__4087 (
            .O(N__16991),
            .I(Lab_UT_di_Mtens_1));
    LocalMux I__4086 (
            .O(N__16982),
            .I(Lab_UT_di_Mtens_1));
    InMux I__4085 (
            .O(N__16977),
            .I(N__16974));
    LocalMux I__4084 (
            .O(N__16974),
            .I(\Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJZ0Z_0 ));
    InMux I__4083 (
            .O(N__16971),
            .I(N__16967));
    InMux I__4082 (
            .O(N__16970),
            .I(N__16960));
    LocalMux I__4081 (
            .O(N__16967),
            .I(N__16957));
    InMux I__4080 (
            .O(N__16966),
            .I(N__16954));
    CascadeMux I__4079 (
            .O(N__16965),
            .I(N__16950));
    CascadeMux I__4078 (
            .O(N__16964),
            .I(N__16947));
    CascadeMux I__4077 (
            .O(N__16963),
            .I(N__16943));
    LocalMux I__4076 (
            .O(N__16960),
            .I(N__16940));
    Span4Mux_v I__4075 (
            .O(N__16957),
            .I(N__16933));
    LocalMux I__4074 (
            .O(N__16954),
            .I(N__16933));
    InMux I__4073 (
            .O(N__16953),
            .I(N__16917));
    InMux I__4072 (
            .O(N__16950),
            .I(N__16917));
    InMux I__4071 (
            .O(N__16947),
            .I(N__16917));
    InMux I__4070 (
            .O(N__16946),
            .I(N__16917));
    InMux I__4069 (
            .O(N__16943),
            .I(N__16917));
    Span4Mux_v I__4068 (
            .O(N__16940),
            .I(N__16914));
    InMux I__4067 (
            .O(N__16939),
            .I(N__16911));
    InMux I__4066 (
            .O(N__16938),
            .I(N__16908));
    Span4Mux_h I__4065 (
            .O(N__16933),
            .I(N__16905));
    InMux I__4064 (
            .O(N__16932),
            .I(N__16902));
    InMux I__4063 (
            .O(N__16931),
            .I(N__16893));
    InMux I__4062 (
            .O(N__16930),
            .I(N__16893));
    InMux I__4061 (
            .O(N__16929),
            .I(N__16893));
    InMux I__4060 (
            .O(N__16928),
            .I(N__16893));
    LocalMux I__4059 (
            .O(N__16917),
            .I(N__16890));
    Odrv4 I__4058 (
            .O(N__16914),
            .I(Lab_UT_di_Mones_2));
    LocalMux I__4057 (
            .O(N__16911),
            .I(Lab_UT_di_Mones_2));
    LocalMux I__4056 (
            .O(N__16908),
            .I(Lab_UT_di_Mones_2));
    Odrv4 I__4055 (
            .O(N__16905),
            .I(Lab_UT_di_Mones_2));
    LocalMux I__4054 (
            .O(N__16902),
            .I(Lab_UT_di_Mones_2));
    LocalMux I__4053 (
            .O(N__16893),
            .I(Lab_UT_di_Mones_2));
    Odrv4 I__4052 (
            .O(N__16890),
            .I(Lab_UT_di_Mones_2));
    InMux I__4051 (
            .O(N__16875),
            .I(N__16870));
    InMux I__4050 (
            .O(N__16874),
            .I(N__16867));
    CascadeMux I__4049 (
            .O(N__16873),
            .I(N__16856));
    LocalMux I__4048 (
            .O(N__16870),
            .I(N__16852));
    LocalMux I__4047 (
            .O(N__16867),
            .I(N__16849));
    CascadeMux I__4046 (
            .O(N__16866),
            .I(N__16845));
    CascadeMux I__4045 (
            .O(N__16865),
            .I(N__16842));
    CascadeMux I__4044 (
            .O(N__16864),
            .I(N__16837));
    InMux I__4043 (
            .O(N__16863),
            .I(N__16826));
    InMux I__4042 (
            .O(N__16862),
            .I(N__16826));
    InMux I__4041 (
            .O(N__16861),
            .I(N__16826));
    InMux I__4040 (
            .O(N__16860),
            .I(N__16826));
    InMux I__4039 (
            .O(N__16859),
            .I(N__16826));
    InMux I__4038 (
            .O(N__16856),
            .I(N__16821));
    InMux I__4037 (
            .O(N__16855),
            .I(N__16821));
    Span4Mux_v I__4036 (
            .O(N__16852),
            .I(N__16816));
    Span4Mux_v I__4035 (
            .O(N__16849),
            .I(N__16816));
    InMux I__4034 (
            .O(N__16848),
            .I(N__16813));
    InMux I__4033 (
            .O(N__16845),
            .I(N__16802));
    InMux I__4032 (
            .O(N__16842),
            .I(N__16802));
    InMux I__4031 (
            .O(N__16841),
            .I(N__16802));
    InMux I__4030 (
            .O(N__16840),
            .I(N__16802));
    InMux I__4029 (
            .O(N__16837),
            .I(N__16802));
    LocalMux I__4028 (
            .O(N__16826),
            .I(N__16799));
    LocalMux I__4027 (
            .O(N__16821),
            .I(Lab_UT_di_Mones_1));
    Odrv4 I__4026 (
            .O(N__16816),
            .I(Lab_UT_di_Mones_1));
    LocalMux I__4025 (
            .O(N__16813),
            .I(Lab_UT_di_Mones_1));
    LocalMux I__4024 (
            .O(N__16802),
            .I(Lab_UT_di_Mones_1));
    Odrv4 I__4023 (
            .O(N__16799),
            .I(Lab_UT_di_Mones_1));
    CascadeMux I__4022 (
            .O(N__16788),
            .I(N__16785));
    InMux I__4021 (
            .O(N__16785),
            .I(N__16777));
    CascadeMux I__4020 (
            .O(N__16784),
            .I(N__16774));
    CascadeMux I__4019 (
            .O(N__16783),
            .I(N__16771));
    CascadeMux I__4018 (
            .O(N__16782),
            .I(N__16768));
    CascadeMux I__4017 (
            .O(N__16781),
            .I(N__16764));
    InMux I__4016 (
            .O(N__16780),
            .I(N__16761));
    LocalMux I__4015 (
            .O(N__16777),
            .I(N__16758));
    InMux I__4014 (
            .O(N__16774),
            .I(N__16755));
    InMux I__4013 (
            .O(N__16771),
            .I(N__16751));
    InMux I__4012 (
            .O(N__16768),
            .I(N__16744));
    InMux I__4011 (
            .O(N__16767),
            .I(N__16744));
    InMux I__4010 (
            .O(N__16764),
            .I(N__16744));
    LocalMux I__4009 (
            .O(N__16761),
            .I(N__16738));
    Span4Mux_v I__4008 (
            .O(N__16758),
            .I(N__16733));
    LocalMux I__4007 (
            .O(N__16755),
            .I(N__16733));
    InMux I__4006 (
            .O(N__16754),
            .I(N__16730));
    LocalMux I__4005 (
            .O(N__16751),
            .I(N__16725));
    LocalMux I__4004 (
            .O(N__16744),
            .I(N__16725));
    CascadeMux I__4003 (
            .O(N__16743),
            .I(N__16722));
    CascadeMux I__4002 (
            .O(N__16742),
            .I(N__16717));
    InMux I__4001 (
            .O(N__16741),
            .I(N__16713));
    Span4Mux_v I__4000 (
            .O(N__16738),
            .I(N__16708));
    Span4Mux_v I__3999 (
            .O(N__16733),
            .I(N__16708));
    LocalMux I__3998 (
            .O(N__16730),
            .I(N__16703));
    Span4Mux_h I__3997 (
            .O(N__16725),
            .I(N__16703));
    InMux I__3996 (
            .O(N__16722),
            .I(N__16692));
    InMux I__3995 (
            .O(N__16721),
            .I(N__16692));
    InMux I__3994 (
            .O(N__16720),
            .I(N__16692));
    InMux I__3993 (
            .O(N__16717),
            .I(N__16692));
    InMux I__3992 (
            .O(N__16716),
            .I(N__16692));
    LocalMux I__3991 (
            .O(N__16713),
            .I(Lab_UT_di_Mones_3));
    Odrv4 I__3990 (
            .O(N__16708),
            .I(Lab_UT_di_Mones_3));
    Odrv4 I__3989 (
            .O(N__16703),
            .I(Lab_UT_di_Mones_3));
    LocalMux I__3988 (
            .O(N__16692),
            .I(Lab_UT_di_Mones_3));
    InMux I__3987 (
            .O(N__16683),
            .I(N__16678));
    InMux I__3986 (
            .O(N__16682),
            .I(N__16675));
    CascadeMux I__3985 (
            .O(N__16681),
            .I(N__16665));
    LocalMux I__3984 (
            .O(N__16678),
            .I(N__16662));
    LocalMux I__3983 (
            .O(N__16675),
            .I(N__16653));
    InMux I__3982 (
            .O(N__16674),
            .I(N__16642));
    InMux I__3981 (
            .O(N__16673),
            .I(N__16642));
    InMux I__3980 (
            .O(N__16672),
            .I(N__16642));
    InMux I__3979 (
            .O(N__16671),
            .I(N__16642));
    InMux I__3978 (
            .O(N__16670),
            .I(N__16642));
    InMux I__3977 (
            .O(N__16669),
            .I(N__16639));
    InMux I__3976 (
            .O(N__16668),
            .I(N__16636));
    InMux I__3975 (
            .O(N__16665),
            .I(N__16633));
    Span4Mux_h I__3974 (
            .O(N__16662),
            .I(N__16630));
    InMux I__3973 (
            .O(N__16661),
            .I(N__16627));
    InMux I__3972 (
            .O(N__16660),
            .I(N__16616));
    InMux I__3971 (
            .O(N__16659),
            .I(N__16616));
    InMux I__3970 (
            .O(N__16658),
            .I(N__16616));
    InMux I__3969 (
            .O(N__16657),
            .I(N__16616));
    InMux I__3968 (
            .O(N__16656),
            .I(N__16616));
    Span4Mux_h I__3967 (
            .O(N__16653),
            .I(N__16611));
    LocalMux I__3966 (
            .O(N__16642),
            .I(N__16611));
    LocalMux I__3965 (
            .O(N__16639),
            .I(Lab_UT_di_Mones_0));
    LocalMux I__3964 (
            .O(N__16636),
            .I(Lab_UT_di_Mones_0));
    LocalMux I__3963 (
            .O(N__16633),
            .I(Lab_UT_di_Mones_0));
    Odrv4 I__3962 (
            .O(N__16630),
            .I(Lab_UT_di_Mones_0));
    LocalMux I__3961 (
            .O(N__16627),
            .I(Lab_UT_di_Mones_0));
    LocalMux I__3960 (
            .O(N__16616),
            .I(Lab_UT_di_Mones_0));
    Odrv4 I__3959 (
            .O(N__16611),
            .I(Lab_UT_di_Mones_0));
    InMux I__3958 (
            .O(N__16596),
            .I(N__16590));
    InMux I__3957 (
            .O(N__16595),
            .I(N__16590));
    LocalMux I__3956 (
            .O(N__16590),
            .I(N__16587));
    Span12Mux_s3_h I__3955 (
            .O(N__16587),
            .I(N__16584));
    Odrv12 I__3954 (
            .O(N__16584),
            .I(\uu2.N_2160_1_0_0 ));
    InMux I__3953 (
            .O(N__16581),
            .I(N__16578));
    LocalMux I__3952 (
            .O(N__16578),
            .I(N__16574));
    InMux I__3951 (
            .O(N__16577),
            .I(N__16571));
    Span4Mux_v I__3950 (
            .O(N__16574),
            .I(N__16564));
    LocalMux I__3949 (
            .O(N__16571),
            .I(N__16564));
    InMux I__3948 (
            .O(N__16570),
            .I(N__16561));
    InMux I__3947 (
            .O(N__16569),
            .I(N__16558));
    Span4Mux_h I__3946 (
            .O(N__16564),
            .I(N__16553));
    LocalMux I__3945 (
            .O(N__16561),
            .I(N__16553));
    LocalMux I__3944 (
            .O(N__16558),
            .I(Lab_UT_dicRun));
    Odrv4 I__3943 (
            .O(N__16553),
            .I(Lab_UT_dicRun));
    InMux I__3942 (
            .O(N__16548),
            .I(N__16543));
    InMux I__3941 (
            .O(N__16547),
            .I(N__16538));
    InMux I__3940 (
            .O(N__16546),
            .I(N__16534));
    LocalMux I__3939 (
            .O(N__16543),
            .I(N__16531));
    InMux I__3938 (
            .O(N__16542),
            .I(N__16526));
    InMux I__3937 (
            .O(N__16541),
            .I(N__16526));
    LocalMux I__3936 (
            .O(N__16538),
            .I(N__16523));
    InMux I__3935 (
            .O(N__16537),
            .I(N__16520));
    LocalMux I__3934 (
            .O(N__16534),
            .I(N__16517));
    Span4Mux_v I__3933 (
            .O(N__16531),
            .I(N__16512));
    LocalMux I__3932 (
            .O(N__16526),
            .I(N__16512));
    Span4Mux_v I__3931 (
            .O(N__16523),
            .I(N__16509));
    LocalMux I__3930 (
            .O(N__16520),
            .I(Lab_UT_l_oneSecPluse));
    Odrv12 I__3929 (
            .O(N__16517),
            .I(Lab_UT_l_oneSecPluse));
    Odrv4 I__3928 (
            .O(N__16512),
            .I(Lab_UT_l_oneSecPluse));
    Odrv4 I__3927 (
            .O(N__16509),
            .I(Lab_UT_l_oneSecPluse));
    IoInMux I__3926 (
            .O(N__16500),
            .I(N__16497));
    LocalMux I__3925 (
            .O(N__16497),
            .I(N__16494));
    Odrv4 I__3924 (
            .O(N__16494),
            .I(led_c_4));
    InMux I__3923 (
            .O(N__16491),
            .I(N__16488));
    LocalMux I__3922 (
            .O(N__16488),
            .I(\uu2.un1_w_addr_displaying_46_1 ));
    CascadeMux I__3921 (
            .O(N__16485),
            .I(\uu2.un1_w_addr_displaying_46_1_cascade_ ));
    InMux I__3920 (
            .O(N__16482),
            .I(N__16479));
    LocalMux I__3919 (
            .O(N__16479),
            .I(N__16476));
    Odrv4 I__3918 (
            .O(N__16476),
            .I(\uu2.w_addr_displaying_RNI8U3D2Z0Z_0 ));
    InMux I__3917 (
            .O(N__16473),
            .I(N__16469));
    InMux I__3916 (
            .O(N__16472),
            .I(N__16466));
    LocalMux I__3915 (
            .O(N__16469),
            .I(N__16460));
    LocalMux I__3914 (
            .O(N__16466),
            .I(N__16455));
    InMux I__3913 (
            .O(N__16465),
            .I(N__16450));
    InMux I__3912 (
            .O(N__16464),
            .I(N__16450));
    InMux I__3911 (
            .O(N__16463),
            .I(N__16447));
    Span4Mux_h I__3910 (
            .O(N__16460),
            .I(N__16444));
    InMux I__3909 (
            .O(N__16459),
            .I(N__16441));
    InMux I__3908 (
            .O(N__16458),
            .I(N__16438));
    Span4Mux_h I__3907 (
            .O(N__16455),
            .I(N__16433));
    LocalMux I__3906 (
            .O(N__16450),
            .I(N__16433));
    LocalMux I__3905 (
            .O(N__16447),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    Odrv4 I__3904 (
            .O(N__16444),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    LocalMux I__3903 (
            .O(N__16441),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    LocalMux I__3902 (
            .O(N__16438),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    Odrv4 I__3901 (
            .O(N__16433),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    InMux I__3900 (
            .O(N__16422),
            .I(N__16418));
    InMux I__3899 (
            .O(N__16421),
            .I(N__16410));
    LocalMux I__3898 (
            .O(N__16418),
            .I(N__16406));
    CascadeMux I__3897 (
            .O(N__16417),
            .I(N__16403));
    InMux I__3896 (
            .O(N__16416),
            .I(N__16398));
    InMux I__3895 (
            .O(N__16415),
            .I(N__16398));
    InMux I__3894 (
            .O(N__16414),
            .I(N__16393));
    InMux I__3893 (
            .O(N__16413),
            .I(N__16393));
    LocalMux I__3892 (
            .O(N__16410),
            .I(N__16390));
    InMux I__3891 (
            .O(N__16409),
            .I(N__16387));
    Span4Mux_h I__3890 (
            .O(N__16406),
            .I(N__16384));
    InMux I__3889 (
            .O(N__16403),
            .I(N__16381));
    LocalMux I__3888 (
            .O(N__16398),
            .I(N__16378));
    LocalMux I__3887 (
            .O(N__16393),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    Odrv4 I__3886 (
            .O(N__16390),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    LocalMux I__3885 (
            .O(N__16387),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    Odrv4 I__3884 (
            .O(N__16384),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    LocalMux I__3883 (
            .O(N__16381),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    Odrv4 I__3882 (
            .O(N__16378),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    InMux I__3881 (
            .O(N__16365),
            .I(N__16360));
    CascadeMux I__3880 (
            .O(N__16364),
            .I(N__16357));
    InMux I__3879 (
            .O(N__16363),
            .I(N__16354));
    LocalMux I__3878 (
            .O(N__16360),
            .I(N__16351));
    InMux I__3877 (
            .O(N__16357),
            .I(N__16348));
    LocalMux I__3876 (
            .O(N__16354),
            .I(N__16337));
    Span4Mux_h I__3875 (
            .O(N__16351),
            .I(N__16337));
    LocalMux I__3874 (
            .O(N__16348),
            .I(N__16334));
    InMux I__3873 (
            .O(N__16347),
            .I(N__16329));
    InMux I__3872 (
            .O(N__16346),
            .I(N__16329));
    InMux I__3871 (
            .O(N__16345),
            .I(N__16320));
    InMux I__3870 (
            .O(N__16344),
            .I(N__16320));
    InMux I__3869 (
            .O(N__16343),
            .I(N__16320));
    InMux I__3868 (
            .O(N__16342),
            .I(N__16320));
    Odrv4 I__3867 (
            .O(N__16337),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    Odrv4 I__3866 (
            .O(N__16334),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__3865 (
            .O(N__16329),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__3864 (
            .O(N__16320),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    InMux I__3863 (
            .O(N__16311),
            .I(N__16308));
    LocalMux I__3862 (
            .O(N__16308),
            .I(\uu2.un1_w_addr_displaying_38_1 ));
    InMux I__3861 (
            .O(N__16305),
            .I(N__16302));
    LocalMux I__3860 (
            .O(N__16302),
            .I(N__16299));
    Span4Mux_v I__3859 (
            .O(N__16299),
            .I(N__16296));
    Odrv4 I__3858 (
            .O(N__16296),
            .I(\uu2.segment3_m_3Z0Z_1 ));
    CascadeMux I__3857 (
            .O(N__16293),
            .I(\uu2.un1_w_addr_displaying_38_1_cascade_ ));
    InMux I__3856 (
            .O(N__16290),
            .I(N__16280));
    InMux I__3855 (
            .O(N__16289),
            .I(N__16269));
    InMux I__3854 (
            .O(N__16288),
            .I(N__16269));
    InMux I__3853 (
            .O(N__16287),
            .I(N__16269));
    InMux I__3852 (
            .O(N__16286),
            .I(N__16269));
    InMux I__3851 (
            .O(N__16285),
            .I(N__16262));
    InMux I__3850 (
            .O(N__16284),
            .I(N__16262));
    InMux I__3849 (
            .O(N__16283),
            .I(N__16262));
    LocalMux I__3848 (
            .O(N__16280),
            .I(N__16259));
    InMux I__3847 (
            .O(N__16279),
            .I(N__16254));
    InMux I__3846 (
            .O(N__16278),
            .I(N__16254));
    LocalMux I__3845 (
            .O(N__16269),
            .I(N__16248));
    LocalMux I__3844 (
            .O(N__16262),
            .I(N__16245));
    Span4Mux_h I__3843 (
            .O(N__16259),
            .I(N__16240));
    LocalMux I__3842 (
            .O(N__16254),
            .I(N__16240));
    InMux I__3841 (
            .O(N__16253),
            .I(N__16237));
    InMux I__3840 (
            .O(N__16252),
            .I(N__16234));
    InMux I__3839 (
            .O(N__16251),
            .I(N__16231));
    Span4Mux_h I__3838 (
            .O(N__16248),
            .I(N__16228));
    Span4Mux_v I__3837 (
            .O(N__16245),
            .I(N__16225));
    Span4Mux_h I__3836 (
            .O(N__16240),
            .I(N__16218));
    LocalMux I__3835 (
            .O(N__16237),
            .I(N__16218));
    LocalMux I__3834 (
            .O(N__16234),
            .I(N__16218));
    LocalMux I__3833 (
            .O(N__16231),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3832 (
            .O(N__16228),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3831 (
            .O(N__16225),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3830 (
            .O(N__16218),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    InMux I__3829 (
            .O(N__16209),
            .I(N__16206));
    LocalMux I__3828 (
            .O(N__16206),
            .I(\uu2.segment3_m_1 ));
    InMux I__3827 (
            .O(N__16203),
            .I(N__16194));
    InMux I__3826 (
            .O(N__16202),
            .I(N__16194));
    InMux I__3825 (
            .O(N__16201),
            .I(N__16188));
    InMux I__3824 (
            .O(N__16200),
            .I(N__16188));
    CascadeMux I__3823 (
            .O(N__16199),
            .I(N__16185));
    LocalMux I__3822 (
            .O(N__16194),
            .I(N__16180));
    InMux I__3821 (
            .O(N__16193),
            .I(N__16177));
    LocalMux I__3820 (
            .O(N__16188),
            .I(N__16172));
    InMux I__3819 (
            .O(N__16185),
            .I(N__16167));
    InMux I__3818 (
            .O(N__16184),
            .I(N__16167));
    InMux I__3817 (
            .O(N__16183),
            .I(N__16164));
    Span4Mux_h I__3816 (
            .O(N__16180),
            .I(N__16161));
    LocalMux I__3815 (
            .O(N__16177),
            .I(N__16158));
    InMux I__3814 (
            .O(N__16176),
            .I(N__16153));
    InMux I__3813 (
            .O(N__16175),
            .I(N__16153));
    Span4Mux_v I__3812 (
            .O(N__16172),
            .I(N__16147));
    LocalMux I__3811 (
            .O(N__16167),
            .I(N__16147));
    LocalMux I__3810 (
            .O(N__16164),
            .I(N__16144));
    Span4Mux_v I__3809 (
            .O(N__16161),
            .I(N__16137));
    Span4Mux_h I__3808 (
            .O(N__16158),
            .I(N__16137));
    LocalMux I__3807 (
            .O(N__16153),
            .I(N__16137));
    InMux I__3806 (
            .O(N__16152),
            .I(N__16131));
    Span4Mux_h I__3805 (
            .O(N__16147),
            .I(N__16128));
    Span12Mux_s11_v I__3804 (
            .O(N__16144),
            .I(N__16125));
    Span4Mux_h I__3803 (
            .O(N__16137),
            .I(N__16122));
    InMux I__3802 (
            .O(N__16136),
            .I(N__16115));
    InMux I__3801 (
            .O(N__16135),
            .I(N__16115));
    InMux I__3800 (
            .O(N__16134),
            .I(N__16115));
    LocalMux I__3799 (
            .O(N__16131),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__3798 (
            .O(N__16128),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv12 I__3797 (
            .O(N__16125),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__3796 (
            .O(N__16122),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__3795 (
            .O(N__16115),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    CascadeMux I__3794 (
            .O(N__16104),
            .I(N__16099));
    InMux I__3793 (
            .O(N__16103),
            .I(N__16087));
    InMux I__3792 (
            .O(N__16102),
            .I(N__16084));
    InMux I__3791 (
            .O(N__16099),
            .I(N__16079));
    InMux I__3790 (
            .O(N__16098),
            .I(N__16076));
    CascadeMux I__3789 (
            .O(N__16097),
            .I(N__16073));
    CascadeMux I__3788 (
            .O(N__16096),
            .I(N__16070));
    CascadeMux I__3787 (
            .O(N__16095),
            .I(N__16067));
    InMux I__3786 (
            .O(N__16094),
            .I(N__16060));
    InMux I__3785 (
            .O(N__16093),
            .I(N__16060));
    CascadeMux I__3784 (
            .O(N__16092),
            .I(N__16050));
    CascadeMux I__3783 (
            .O(N__16091),
            .I(N__16046));
    InMux I__3782 (
            .O(N__16090),
            .I(N__16042));
    LocalMux I__3781 (
            .O(N__16087),
            .I(N__16037));
    LocalMux I__3780 (
            .O(N__16084),
            .I(N__16037));
    InMux I__3779 (
            .O(N__16083),
            .I(N__16032));
    InMux I__3778 (
            .O(N__16082),
            .I(N__16032));
    LocalMux I__3777 (
            .O(N__16079),
            .I(N__16029));
    LocalMux I__3776 (
            .O(N__16076),
            .I(N__16026));
    InMux I__3775 (
            .O(N__16073),
            .I(N__16023));
    InMux I__3774 (
            .O(N__16070),
            .I(N__16014));
    InMux I__3773 (
            .O(N__16067),
            .I(N__16014));
    InMux I__3772 (
            .O(N__16066),
            .I(N__16014));
    InMux I__3771 (
            .O(N__16065),
            .I(N__16014));
    LocalMux I__3770 (
            .O(N__16060),
            .I(N__16011));
    InMux I__3769 (
            .O(N__16059),
            .I(N__16006));
    InMux I__3768 (
            .O(N__16058),
            .I(N__16006));
    InMux I__3767 (
            .O(N__16057),
            .I(N__16001));
    InMux I__3766 (
            .O(N__16056),
            .I(N__16001));
    InMux I__3765 (
            .O(N__16055),
            .I(N__15994));
    InMux I__3764 (
            .O(N__16054),
            .I(N__15994));
    InMux I__3763 (
            .O(N__16053),
            .I(N__15994));
    InMux I__3762 (
            .O(N__16050),
            .I(N__15989));
    InMux I__3761 (
            .O(N__16049),
            .I(N__15989));
    InMux I__3760 (
            .O(N__16046),
            .I(N__15984));
    InMux I__3759 (
            .O(N__16045),
            .I(N__15984));
    LocalMux I__3758 (
            .O(N__16042),
            .I(N__15981));
    Span4Mux_v I__3757 (
            .O(N__16037),
            .I(N__15978));
    LocalMux I__3756 (
            .O(N__16032),
            .I(N__15971));
    Span4Mux_v I__3755 (
            .O(N__16029),
            .I(N__15971));
    Span4Mux_h I__3754 (
            .O(N__16026),
            .I(N__15971));
    LocalMux I__3753 (
            .O(N__16023),
            .I(N__15964));
    LocalMux I__3752 (
            .O(N__16014),
            .I(N__15964));
    Span4Mux_v I__3751 (
            .O(N__16011),
            .I(N__15964));
    LocalMux I__3750 (
            .O(N__16006),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__3749 (
            .O(N__16001),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__3748 (
            .O(N__15994),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__3747 (
            .O(N__15989),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__3746 (
            .O(N__15984),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__3745 (
            .O(N__15981),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__3744 (
            .O(N__15978),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__3743 (
            .O(N__15971),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__3742 (
            .O(N__15964),
            .I(\uu2.un21_w_addr_displaying_i ));
    InMux I__3741 (
            .O(N__15945),
            .I(N__15940));
    InMux I__3740 (
            .O(N__15944),
            .I(N__15937));
    InMux I__3739 (
            .O(N__15943),
            .I(N__15934));
    LocalMux I__3738 (
            .O(N__15940),
            .I(N__15931));
    LocalMux I__3737 (
            .O(N__15937),
            .I(N__15928));
    LocalMux I__3736 (
            .O(N__15934),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    Odrv4 I__3735 (
            .O(N__15931),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    Odrv4 I__3734 (
            .O(N__15928),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    InMux I__3733 (
            .O(N__15921),
            .I(N__15914));
    InMux I__3732 (
            .O(N__15920),
            .I(N__15911));
    InMux I__3731 (
            .O(N__15919),
            .I(N__15906));
    InMux I__3730 (
            .O(N__15918),
            .I(N__15906));
    InMux I__3729 (
            .O(N__15917),
            .I(N__15903));
    LocalMux I__3728 (
            .O(N__15914),
            .I(N__15869));
    LocalMux I__3727 (
            .O(N__15911),
            .I(N__15866));
    LocalMux I__3726 (
            .O(N__15906),
            .I(N__15863));
    LocalMux I__3725 (
            .O(N__15903),
            .I(N__15860));
    SRMux I__3724 (
            .O(N__15902),
            .I(N__15753));
    SRMux I__3723 (
            .O(N__15901),
            .I(N__15753));
    SRMux I__3722 (
            .O(N__15900),
            .I(N__15753));
    SRMux I__3721 (
            .O(N__15899),
            .I(N__15753));
    SRMux I__3720 (
            .O(N__15898),
            .I(N__15753));
    SRMux I__3719 (
            .O(N__15897),
            .I(N__15753));
    SRMux I__3718 (
            .O(N__15896),
            .I(N__15753));
    SRMux I__3717 (
            .O(N__15895),
            .I(N__15753));
    SRMux I__3716 (
            .O(N__15894),
            .I(N__15753));
    SRMux I__3715 (
            .O(N__15893),
            .I(N__15753));
    SRMux I__3714 (
            .O(N__15892),
            .I(N__15753));
    SRMux I__3713 (
            .O(N__15891),
            .I(N__15753));
    SRMux I__3712 (
            .O(N__15890),
            .I(N__15753));
    SRMux I__3711 (
            .O(N__15889),
            .I(N__15753));
    SRMux I__3710 (
            .O(N__15888),
            .I(N__15753));
    SRMux I__3709 (
            .O(N__15887),
            .I(N__15753));
    SRMux I__3708 (
            .O(N__15886),
            .I(N__15753));
    SRMux I__3707 (
            .O(N__15885),
            .I(N__15753));
    SRMux I__3706 (
            .O(N__15884),
            .I(N__15753));
    SRMux I__3705 (
            .O(N__15883),
            .I(N__15753));
    SRMux I__3704 (
            .O(N__15882),
            .I(N__15753));
    SRMux I__3703 (
            .O(N__15881),
            .I(N__15753));
    SRMux I__3702 (
            .O(N__15880),
            .I(N__15753));
    SRMux I__3701 (
            .O(N__15879),
            .I(N__15753));
    SRMux I__3700 (
            .O(N__15878),
            .I(N__15753));
    SRMux I__3699 (
            .O(N__15877),
            .I(N__15753));
    SRMux I__3698 (
            .O(N__15876),
            .I(N__15753));
    SRMux I__3697 (
            .O(N__15875),
            .I(N__15753));
    SRMux I__3696 (
            .O(N__15874),
            .I(N__15753));
    SRMux I__3695 (
            .O(N__15873),
            .I(N__15753));
    SRMux I__3694 (
            .O(N__15872),
            .I(N__15753));
    Glb2LocalMux I__3693 (
            .O(N__15869),
            .I(N__15753));
    Glb2LocalMux I__3692 (
            .O(N__15866),
            .I(N__15753));
    Glb2LocalMux I__3691 (
            .O(N__15863),
            .I(N__15753));
    Glb2LocalMux I__3690 (
            .O(N__15860),
            .I(N__15753));
    SRMux I__3689 (
            .O(N__15859),
            .I(N__15753));
    SRMux I__3688 (
            .O(N__15858),
            .I(N__15753));
    SRMux I__3687 (
            .O(N__15857),
            .I(N__15753));
    SRMux I__3686 (
            .O(N__15856),
            .I(N__15753));
    SRMux I__3685 (
            .O(N__15855),
            .I(N__15753));
    SRMux I__3684 (
            .O(N__15854),
            .I(N__15753));
    SRMux I__3683 (
            .O(N__15853),
            .I(N__15753));
    SRMux I__3682 (
            .O(N__15852),
            .I(N__15753));
    SRMux I__3681 (
            .O(N__15851),
            .I(N__15753));
    SRMux I__3680 (
            .O(N__15850),
            .I(N__15753));
    SRMux I__3679 (
            .O(N__15849),
            .I(N__15753));
    SRMux I__3678 (
            .O(N__15848),
            .I(N__15753));
    GlobalMux I__3677 (
            .O(N__15753),
            .I(N__15750));
    gio2CtrlBuf I__3676 (
            .O(N__15750),
            .I(rst_g));
    InMux I__3675 (
            .O(N__15747),
            .I(N__15744));
    LocalMux I__3674 (
            .O(N__15744),
            .I(N__15741));
    Span4Mux_h I__3673 (
            .O(N__15741),
            .I(N__15738));
    Odrv4 I__3672 (
            .O(N__15738),
            .I(\uu2.mem0.N_2160_2 ));
    InMux I__3671 (
            .O(N__15735),
            .I(N__15726));
    InMux I__3670 (
            .O(N__15734),
            .I(N__15716));
    InMux I__3669 (
            .O(N__15733),
            .I(N__15716));
    InMux I__3668 (
            .O(N__15732),
            .I(N__15716));
    InMux I__3667 (
            .O(N__15731),
            .I(N__15716));
    InMux I__3666 (
            .O(N__15730),
            .I(N__15708));
    InMux I__3665 (
            .O(N__15729),
            .I(N__15708));
    LocalMux I__3664 (
            .O(N__15726),
            .I(N__15705));
    InMux I__3663 (
            .O(N__15725),
            .I(N__15702));
    LocalMux I__3662 (
            .O(N__15716),
            .I(N__15699));
    InMux I__3661 (
            .O(N__15715),
            .I(N__15692));
    InMux I__3660 (
            .O(N__15714),
            .I(N__15692));
    InMux I__3659 (
            .O(N__15713),
            .I(N__15692));
    LocalMux I__3658 (
            .O(N__15708),
            .I(N__15686));
    Span4Mux_v I__3657 (
            .O(N__15705),
            .I(N__15681));
    LocalMux I__3656 (
            .O(N__15702),
            .I(N__15681));
    Span12Mux_s9_v I__3655 (
            .O(N__15699),
            .I(N__15678));
    LocalMux I__3654 (
            .O(N__15692),
            .I(N__15675));
    InMux I__3653 (
            .O(N__15691),
            .I(N__15668));
    InMux I__3652 (
            .O(N__15690),
            .I(N__15668));
    InMux I__3651 (
            .O(N__15689),
            .I(N__15668));
    Span4Mux_h I__3650 (
            .O(N__15686),
            .I(N__15665));
    Odrv4 I__3649 (
            .O(N__15681),
            .I(Lab_UT_di_Sones_0));
    Odrv12 I__3648 (
            .O(N__15678),
            .I(Lab_UT_di_Sones_0));
    Odrv12 I__3647 (
            .O(N__15675),
            .I(Lab_UT_di_Sones_0));
    LocalMux I__3646 (
            .O(N__15668),
            .I(Lab_UT_di_Sones_0));
    Odrv4 I__3645 (
            .O(N__15665),
            .I(Lab_UT_di_Sones_0));
    InMux I__3644 (
            .O(N__15654),
            .I(N__15650));
    InMux I__3643 (
            .O(N__15653),
            .I(N__15647));
    LocalMux I__3642 (
            .O(N__15650),
            .I(N__15643));
    LocalMux I__3641 (
            .O(N__15647),
            .I(N__15632));
    InMux I__3640 (
            .O(N__15646),
            .I(N__15629));
    Span4Mux_h I__3639 (
            .O(N__15643),
            .I(N__15623));
    InMux I__3638 (
            .O(N__15642),
            .I(N__15620));
    InMux I__3637 (
            .O(N__15641),
            .I(N__15611));
    InMux I__3636 (
            .O(N__15640),
            .I(N__15611));
    InMux I__3635 (
            .O(N__15639),
            .I(N__15611));
    InMux I__3634 (
            .O(N__15638),
            .I(N__15611));
    InMux I__3633 (
            .O(N__15637),
            .I(N__15603));
    InMux I__3632 (
            .O(N__15636),
            .I(N__15603));
    InMux I__3631 (
            .O(N__15635),
            .I(N__15603));
    Span4Mux_v I__3630 (
            .O(N__15632),
            .I(N__15598));
    LocalMux I__3629 (
            .O(N__15629),
            .I(N__15598));
    InMux I__3628 (
            .O(N__15628),
            .I(N__15591));
    InMux I__3627 (
            .O(N__15627),
            .I(N__15591));
    InMux I__3626 (
            .O(N__15626),
            .I(N__15591));
    Sp12to4 I__3625 (
            .O(N__15623),
            .I(N__15584));
    LocalMux I__3624 (
            .O(N__15620),
            .I(N__15584));
    LocalMux I__3623 (
            .O(N__15611),
            .I(N__15584));
    InMux I__3622 (
            .O(N__15610),
            .I(N__15581));
    LocalMux I__3621 (
            .O(N__15603),
            .I(Lab_UT_di_Stens_0));
    Odrv4 I__3620 (
            .O(N__15598),
            .I(Lab_UT_di_Stens_0));
    LocalMux I__3619 (
            .O(N__15591),
            .I(Lab_UT_di_Stens_0));
    Odrv12 I__3618 (
            .O(N__15584),
            .I(Lab_UT_di_Stens_0));
    LocalMux I__3617 (
            .O(N__15581),
            .I(Lab_UT_di_Stens_0));
    InMux I__3616 (
            .O(N__15570),
            .I(N__15567));
    LocalMux I__3615 (
            .O(N__15567),
            .I(\uu2.w_addr_displaying_4_rep2_RNI4S6JZ0 ));
    CascadeMux I__3614 (
            .O(N__15564),
            .I(\uu2.w_addr_displaying_fast_RNIEDBMZ0Z_7_cascade_ ));
    InMux I__3613 (
            .O(N__15561),
            .I(N__15558));
    LocalMux I__3612 (
            .O(N__15558),
            .I(N__15555));
    Odrv4 I__3611 (
            .O(N__15555),
            .I(\uu2.un1_segment4_sn_N_38_0 ));
    CascadeMux I__3610 (
            .O(N__15552),
            .I(N__15548));
    InMux I__3609 (
            .O(N__15551),
            .I(N__15540));
    InMux I__3608 (
            .O(N__15548),
            .I(N__15540));
    InMux I__3607 (
            .O(N__15547),
            .I(N__15537));
    CascadeMux I__3606 (
            .O(N__15546),
            .I(N__15534));
    CascadeMux I__3605 (
            .O(N__15545),
            .I(N__15527));
    LocalMux I__3604 (
            .O(N__15540),
            .I(N__15523));
    LocalMux I__3603 (
            .O(N__15537),
            .I(N__15520));
    InMux I__3602 (
            .O(N__15534),
            .I(N__15515));
    InMux I__3601 (
            .O(N__15533),
            .I(N__15515));
    InMux I__3600 (
            .O(N__15532),
            .I(N__15510));
    InMux I__3599 (
            .O(N__15531),
            .I(N__15510));
    InMux I__3598 (
            .O(N__15530),
            .I(N__15503));
    InMux I__3597 (
            .O(N__15527),
            .I(N__15503));
    InMux I__3596 (
            .O(N__15526),
            .I(N__15503));
    Odrv4 I__3595 (
            .O(N__15523),
            .I(\uu2.w_addr_displaying_4_repZ0Z2 ));
    Odrv4 I__3594 (
            .O(N__15520),
            .I(\uu2.w_addr_displaying_4_repZ0Z2 ));
    LocalMux I__3593 (
            .O(N__15515),
            .I(\uu2.w_addr_displaying_4_repZ0Z2 ));
    LocalMux I__3592 (
            .O(N__15510),
            .I(\uu2.w_addr_displaying_4_repZ0Z2 ));
    LocalMux I__3591 (
            .O(N__15503),
            .I(\uu2.w_addr_displaying_4_repZ0Z2 ));
    InMux I__3590 (
            .O(N__15492),
            .I(N__15487));
    InMux I__3589 (
            .O(N__15491),
            .I(N__15484));
    CascadeMux I__3588 (
            .O(N__15490),
            .I(N__15481));
    LocalMux I__3587 (
            .O(N__15487),
            .I(N__15477));
    LocalMux I__3586 (
            .O(N__15484),
            .I(N__15474));
    InMux I__3585 (
            .O(N__15481),
            .I(N__15471));
    InMux I__3584 (
            .O(N__15480),
            .I(N__15468));
    Odrv4 I__3583 (
            .O(N__15477),
            .I(\uu2.N_111 ));
    Odrv4 I__3582 (
            .O(N__15474),
            .I(\uu2.N_111 ));
    LocalMux I__3581 (
            .O(N__15471),
            .I(\uu2.N_111 ));
    LocalMux I__3580 (
            .O(N__15468),
            .I(\uu2.N_111 ));
    InMux I__3579 (
            .O(N__15459),
            .I(N__15453));
    InMux I__3578 (
            .O(N__15458),
            .I(N__15446));
    InMux I__3577 (
            .O(N__15457),
            .I(N__15443));
    CascadeMux I__3576 (
            .O(N__15456),
            .I(N__15438));
    LocalMux I__3575 (
            .O(N__15453),
            .I(N__15435));
    InMux I__3574 (
            .O(N__15452),
            .I(N__15432));
    InMux I__3573 (
            .O(N__15451),
            .I(N__15427));
    InMux I__3572 (
            .O(N__15450),
            .I(N__15427));
    CascadeMux I__3571 (
            .O(N__15449),
            .I(N__15422));
    LocalMux I__3570 (
            .O(N__15446),
            .I(N__15415));
    LocalMux I__3569 (
            .O(N__15443),
            .I(N__15415));
    InMux I__3568 (
            .O(N__15442),
            .I(N__15412));
    InMux I__3567 (
            .O(N__15441),
            .I(N__15409));
    InMux I__3566 (
            .O(N__15438),
            .I(N__15406));
    Span4Mux_h I__3565 (
            .O(N__15435),
            .I(N__15403));
    LocalMux I__3564 (
            .O(N__15432),
            .I(N__15398));
    LocalMux I__3563 (
            .O(N__15427),
            .I(N__15398));
    InMux I__3562 (
            .O(N__15426),
            .I(N__15393));
    InMux I__3561 (
            .O(N__15425),
            .I(N__15393));
    InMux I__3560 (
            .O(N__15422),
            .I(N__15386));
    InMux I__3559 (
            .O(N__15421),
            .I(N__15386));
    InMux I__3558 (
            .O(N__15420),
            .I(N__15386));
    Odrv4 I__3557 (
            .O(N__15415),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__3556 (
            .O(N__15412),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__3555 (
            .O(N__15409),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__3554 (
            .O(N__15406),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__3553 (
            .O(N__15403),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__3552 (
            .O(N__15398),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__3551 (
            .O(N__15393),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__3550 (
            .O(N__15386),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    InMux I__3549 (
            .O(N__15369),
            .I(N__15362));
    CascadeMux I__3548 (
            .O(N__15368),
            .I(N__15359));
    InMux I__3547 (
            .O(N__15367),
            .I(N__15356));
    InMux I__3546 (
            .O(N__15366),
            .I(N__15353));
    InMux I__3545 (
            .O(N__15365),
            .I(N__15350));
    LocalMux I__3544 (
            .O(N__15362),
            .I(N__15347));
    InMux I__3543 (
            .O(N__15359),
            .I(N__15342));
    LocalMux I__3542 (
            .O(N__15356),
            .I(N__15339));
    LocalMux I__3541 (
            .O(N__15353),
            .I(N__15334));
    LocalMux I__3540 (
            .O(N__15350),
            .I(N__15334));
    Span4Mux_v I__3539 (
            .O(N__15347),
            .I(N__15331));
    InMux I__3538 (
            .O(N__15346),
            .I(N__15326));
    InMux I__3537 (
            .O(N__15345),
            .I(N__15326));
    LocalMux I__3536 (
            .O(N__15342),
            .I(N__15321));
    Span4Mux_h I__3535 (
            .O(N__15339),
            .I(N__15321));
    Span4Mux_v I__3534 (
            .O(N__15334),
            .I(N__15318));
    Odrv4 I__3533 (
            .O(N__15331),
            .I(\uu2.Z_decfrac106_6 ));
    LocalMux I__3532 (
            .O(N__15326),
            .I(\uu2.Z_decfrac106_6 ));
    Odrv4 I__3531 (
            .O(N__15321),
            .I(\uu2.Z_decfrac106_6 ));
    Odrv4 I__3530 (
            .O(N__15318),
            .I(\uu2.Z_decfrac106_6 ));
    CascadeMux I__3529 (
            .O(N__15309),
            .I(N__15302));
    InMux I__3528 (
            .O(N__15308),
            .I(N__15296));
    InMux I__3527 (
            .O(N__15307),
            .I(N__15296));
    CascadeMux I__3526 (
            .O(N__15306),
            .I(N__15293));
    InMux I__3525 (
            .O(N__15305),
            .I(N__15288));
    InMux I__3524 (
            .O(N__15302),
            .I(N__15283));
    InMux I__3523 (
            .O(N__15301),
            .I(N__15283));
    LocalMux I__3522 (
            .O(N__15296),
            .I(N__15280));
    InMux I__3521 (
            .O(N__15293),
            .I(N__15275));
    InMux I__3520 (
            .O(N__15292),
            .I(N__15275));
    InMux I__3519 (
            .O(N__15291),
            .I(N__15272));
    LocalMux I__3518 (
            .O(N__15288),
            .I(N__15267));
    LocalMux I__3517 (
            .O(N__15283),
            .I(N__15267));
    Span4Mux_h I__3516 (
            .O(N__15280),
            .I(N__15264));
    LocalMux I__3515 (
            .O(N__15275),
            .I(N__15261));
    LocalMux I__3514 (
            .O(N__15272),
            .I(N__15256));
    Span4Mux_h I__3513 (
            .O(N__15267),
            .I(N__15256));
    Odrv4 I__3512 (
            .O(N__15264),
            .I(\uu2.un15_w_data_displaying_5 ));
    Odrv4 I__3511 (
            .O(N__15261),
            .I(\uu2.un15_w_data_displaying_5 ));
    Odrv4 I__3510 (
            .O(N__15256),
            .I(\uu2.un15_w_data_displaying_5 ));
    InMux I__3509 (
            .O(N__15249),
            .I(N__15244));
    InMux I__3508 (
            .O(N__15248),
            .I(N__15241));
    CascadeMux I__3507 (
            .O(N__15247),
            .I(N__15237));
    LocalMux I__3506 (
            .O(N__15244),
            .I(N__15232));
    LocalMux I__3505 (
            .O(N__15241),
            .I(N__15229));
    CascadeMux I__3504 (
            .O(N__15240),
            .I(N__15226));
    InMux I__3503 (
            .O(N__15237),
            .I(N__15223));
    InMux I__3502 (
            .O(N__15236),
            .I(N__15218));
    InMux I__3501 (
            .O(N__15235),
            .I(N__15218));
    Span4Mux_h I__3500 (
            .O(N__15232),
            .I(N__15215));
    Span4Mux_h I__3499 (
            .O(N__15229),
            .I(N__15212));
    InMux I__3498 (
            .O(N__15226),
            .I(N__15209));
    LocalMux I__3497 (
            .O(N__15223),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    LocalMux I__3496 (
            .O(N__15218),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    Odrv4 I__3495 (
            .O(N__15215),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    Odrv4 I__3494 (
            .O(N__15212),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    LocalMux I__3493 (
            .O(N__15209),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    CascadeMux I__3492 (
            .O(N__15198),
            .I(L3_segment4_2_cascade_));
    InMux I__3491 (
            .O(N__15195),
            .I(N__15192));
    LocalMux I__3490 (
            .O(N__15192),
            .I(\uu2.N_280 ));
    CascadeMux I__3489 (
            .O(N__15189),
            .I(N__15184));
    InMux I__3488 (
            .O(N__15188),
            .I(N__15179));
    InMux I__3487 (
            .O(N__15187),
            .I(N__15176));
    InMux I__3486 (
            .O(N__15184),
            .I(N__15173));
    InMux I__3485 (
            .O(N__15183),
            .I(N__15168));
    InMux I__3484 (
            .O(N__15182),
            .I(N__15168));
    LocalMux I__3483 (
            .O(N__15179),
            .I(N__15163));
    LocalMux I__3482 (
            .O(N__15176),
            .I(N__15160));
    LocalMux I__3481 (
            .O(N__15173),
            .I(N__15157));
    LocalMux I__3480 (
            .O(N__15168),
            .I(N__15154));
    InMux I__3479 (
            .O(N__15167),
            .I(N__15149));
    InMux I__3478 (
            .O(N__15166),
            .I(N__15149));
    Span4Mux_v I__3477 (
            .O(N__15163),
            .I(N__15138));
    Span4Mux_h I__3476 (
            .O(N__15160),
            .I(N__15138));
    Span4Mux_h I__3475 (
            .O(N__15157),
            .I(N__15138));
    Span4Mux_h I__3474 (
            .O(N__15154),
            .I(N__15138));
    LocalMux I__3473 (
            .O(N__15149),
            .I(N__15138));
    Span4Mux_v I__3472 (
            .O(N__15138),
            .I(N__15127));
    InMux I__3471 (
            .O(N__15137),
            .I(N__15120));
    InMux I__3470 (
            .O(N__15136),
            .I(N__15120));
    InMux I__3469 (
            .O(N__15135),
            .I(N__15120));
    InMux I__3468 (
            .O(N__15134),
            .I(N__15109));
    InMux I__3467 (
            .O(N__15133),
            .I(N__15109));
    InMux I__3466 (
            .O(N__15132),
            .I(N__15109));
    InMux I__3465 (
            .O(N__15131),
            .I(N__15109));
    InMux I__3464 (
            .O(N__15130),
            .I(N__15109));
    Odrv4 I__3463 (
            .O(N__15127),
            .I(Lab_UT_di_Mtens_2));
    LocalMux I__3462 (
            .O(N__15120),
            .I(Lab_UT_di_Mtens_2));
    LocalMux I__3461 (
            .O(N__15109),
            .I(Lab_UT_di_Mtens_2));
    CascadeMux I__3460 (
            .O(N__15102),
            .I(N__15096));
    CascadeMux I__3459 (
            .O(N__15101),
            .I(N__15092));
    CascadeMux I__3458 (
            .O(N__15100),
            .I(N__15089));
    InMux I__3457 (
            .O(N__15099),
            .I(N__15085));
    InMux I__3456 (
            .O(N__15096),
            .I(N__15082));
    InMux I__3455 (
            .O(N__15095),
            .I(N__15079));
    InMux I__3454 (
            .O(N__15092),
            .I(N__15074));
    InMux I__3453 (
            .O(N__15089),
            .I(N__15074));
    CascadeMux I__3452 (
            .O(N__15088),
            .I(N__15070));
    LocalMux I__3451 (
            .O(N__15085),
            .I(N__15067));
    LocalMux I__3450 (
            .O(N__15082),
            .I(N__15064));
    LocalMux I__3449 (
            .O(N__15079),
            .I(N__15061));
    LocalMux I__3448 (
            .O(N__15074),
            .I(N__15058));
    InMux I__3447 (
            .O(N__15073),
            .I(N__15053));
    InMux I__3446 (
            .O(N__15070),
            .I(N__15053));
    Span4Mux_v I__3445 (
            .O(N__15067),
            .I(N__15043));
    Span4Mux_h I__3444 (
            .O(N__15064),
            .I(N__15034));
    Span4Mux_h I__3443 (
            .O(N__15061),
            .I(N__15034));
    Span4Mux_h I__3442 (
            .O(N__15058),
            .I(N__15034));
    LocalMux I__3441 (
            .O(N__15053),
            .I(N__15034));
    InMux I__3440 (
            .O(N__15052),
            .I(N__15027));
    InMux I__3439 (
            .O(N__15051),
            .I(N__15027));
    InMux I__3438 (
            .O(N__15050),
            .I(N__15027));
    InMux I__3437 (
            .O(N__15049),
            .I(N__15018));
    InMux I__3436 (
            .O(N__15048),
            .I(N__15018));
    InMux I__3435 (
            .O(N__15047),
            .I(N__15018));
    InMux I__3434 (
            .O(N__15046),
            .I(N__15018));
    Odrv4 I__3433 (
            .O(N__15043),
            .I(Lab_UT_di_Mtens_3));
    Odrv4 I__3432 (
            .O(N__15034),
            .I(Lab_UT_di_Mtens_3));
    LocalMux I__3431 (
            .O(N__15027),
            .I(Lab_UT_di_Mtens_3));
    LocalMux I__3430 (
            .O(N__15018),
            .I(Lab_UT_di_Mtens_3));
    InMux I__3429 (
            .O(N__15009),
            .I(N__15006));
    LocalMux I__3428 (
            .O(N__15006),
            .I(L3_segment4_4));
    InMux I__3427 (
            .O(N__15003),
            .I(N__14995));
    CascadeMux I__3426 (
            .O(N__15002),
            .I(N__14989));
    InMux I__3425 (
            .O(N__15001),
            .I(N__14984));
    InMux I__3424 (
            .O(N__15000),
            .I(N__14979));
    InMux I__3423 (
            .O(N__14999),
            .I(N__14979));
    InMux I__3422 (
            .O(N__14998),
            .I(N__14976));
    LocalMux I__3421 (
            .O(N__14995),
            .I(N__14972));
    InMux I__3420 (
            .O(N__14994),
            .I(N__14965));
    InMux I__3419 (
            .O(N__14993),
            .I(N__14965));
    InMux I__3418 (
            .O(N__14992),
            .I(N__14965));
    InMux I__3417 (
            .O(N__14989),
            .I(N__14962));
    InMux I__3416 (
            .O(N__14988),
            .I(N__14958));
    CascadeMux I__3415 (
            .O(N__14987),
            .I(N__14955));
    LocalMux I__3414 (
            .O(N__14984),
            .I(N__14950));
    LocalMux I__3413 (
            .O(N__14979),
            .I(N__14950));
    LocalMux I__3412 (
            .O(N__14976),
            .I(N__14947));
    InMux I__3411 (
            .O(N__14975),
            .I(N__14944));
    Span4Mux_v I__3410 (
            .O(N__14972),
            .I(N__14937));
    LocalMux I__3409 (
            .O(N__14965),
            .I(N__14937));
    LocalMux I__3408 (
            .O(N__14962),
            .I(N__14937));
    InMux I__3407 (
            .O(N__14961),
            .I(N__14934));
    LocalMux I__3406 (
            .O(N__14958),
            .I(N__14931));
    InMux I__3405 (
            .O(N__14955),
            .I(N__14928));
    Span4Mux_h I__3404 (
            .O(N__14950),
            .I(N__14925));
    Span4Mux_h I__3403 (
            .O(N__14947),
            .I(N__14918));
    LocalMux I__3402 (
            .O(N__14944),
            .I(N__14918));
    Span4Mux_h I__3401 (
            .O(N__14937),
            .I(N__14918));
    LocalMux I__3400 (
            .O(N__14934),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__3399 (
            .O(N__14931),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__3398 (
            .O(N__14928),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__3397 (
            .O(N__14925),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__3396 (
            .O(N__14918),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    CascadeMux I__3395 (
            .O(N__14907),
            .I(N__14903));
    InMux I__3394 (
            .O(N__14906),
            .I(N__14897));
    InMux I__3393 (
            .O(N__14903),
            .I(N__14897));
    CascadeMux I__3392 (
            .O(N__14902),
            .I(N__14893));
    LocalMux I__3391 (
            .O(N__14897),
            .I(N__14884));
    InMux I__3390 (
            .O(N__14896),
            .I(N__14881));
    InMux I__3389 (
            .O(N__14893),
            .I(N__14878));
    InMux I__3388 (
            .O(N__14892),
            .I(N__14875));
    InMux I__3387 (
            .O(N__14891),
            .I(N__14870));
    InMux I__3386 (
            .O(N__14890),
            .I(N__14870));
    CascadeMux I__3385 (
            .O(N__14889),
            .I(N__14867));
    InMux I__3384 (
            .O(N__14888),
            .I(N__14861));
    InMux I__3383 (
            .O(N__14887),
            .I(N__14861));
    Span4Mux_v I__3382 (
            .O(N__14884),
            .I(N__14856));
    LocalMux I__3381 (
            .O(N__14881),
            .I(N__14856));
    LocalMux I__3380 (
            .O(N__14878),
            .I(N__14851));
    LocalMux I__3379 (
            .O(N__14875),
            .I(N__14851));
    LocalMux I__3378 (
            .O(N__14870),
            .I(N__14848));
    InMux I__3377 (
            .O(N__14867),
            .I(N__14843));
    InMux I__3376 (
            .O(N__14866),
            .I(N__14843));
    LocalMux I__3375 (
            .O(N__14861),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    Odrv4 I__3374 (
            .O(N__14856),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    Odrv4 I__3373 (
            .O(N__14851),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    Odrv4 I__3372 (
            .O(N__14848),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    LocalMux I__3371 (
            .O(N__14843),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    InMux I__3370 (
            .O(N__14832),
            .I(N__14828));
    CascadeMux I__3369 (
            .O(N__14831),
            .I(N__14823));
    LocalMux I__3368 (
            .O(N__14828),
            .I(N__14817));
    InMux I__3367 (
            .O(N__14827),
            .I(N__14814));
    InMux I__3366 (
            .O(N__14826),
            .I(N__14809));
    InMux I__3365 (
            .O(N__14823),
            .I(N__14809));
    InMux I__3364 (
            .O(N__14822),
            .I(N__14806));
    InMux I__3363 (
            .O(N__14821),
            .I(N__14801));
    InMux I__3362 (
            .O(N__14820),
            .I(N__14801));
    Span4Mux_h I__3361 (
            .O(N__14817),
            .I(N__14796));
    LocalMux I__3360 (
            .O(N__14814),
            .I(N__14796));
    LocalMux I__3359 (
            .O(N__14809),
            .I(N__14793));
    LocalMux I__3358 (
            .O(N__14806),
            .I(N__14787));
    LocalMux I__3357 (
            .O(N__14801),
            .I(N__14780));
    Span4Mux_h I__3356 (
            .O(N__14796),
            .I(N__14780));
    Span4Mux_v I__3355 (
            .O(N__14793),
            .I(N__14780));
    InMux I__3354 (
            .O(N__14792),
            .I(N__14773));
    InMux I__3353 (
            .O(N__14791),
            .I(N__14773));
    InMux I__3352 (
            .O(N__14790),
            .I(N__14773));
    Odrv4 I__3351 (
            .O(N__14787),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    Odrv4 I__3350 (
            .O(N__14780),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    LocalMux I__3349 (
            .O(N__14773),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    CascadeMux I__3348 (
            .O(N__14766),
            .I(N__14763));
    InMux I__3347 (
            .O(N__14763),
            .I(N__14760));
    LocalMux I__3346 (
            .O(N__14760),
            .I(N__14757));
    Span4Mux_h I__3345 (
            .O(N__14757),
            .I(N__14754));
    Odrv4 I__3344 (
            .O(N__14754),
            .I(\uu2.un1_segment3_m4_s_2_1 ));
    InMux I__3343 (
            .O(N__14751),
            .I(N__14738));
    InMux I__3342 (
            .O(N__14750),
            .I(N__14738));
    InMux I__3341 (
            .O(N__14749),
            .I(N__14735));
    InMux I__3340 (
            .O(N__14748),
            .I(N__14721));
    InMux I__3339 (
            .O(N__14747),
            .I(N__14721));
    InMux I__3338 (
            .O(N__14746),
            .I(N__14721));
    InMux I__3337 (
            .O(N__14745),
            .I(N__14721));
    InMux I__3336 (
            .O(N__14744),
            .I(N__14721));
    InMux I__3335 (
            .O(N__14743),
            .I(N__14721));
    LocalMux I__3334 (
            .O(N__14738),
            .I(N__14716));
    LocalMux I__3333 (
            .O(N__14735),
            .I(N__14713));
    InMux I__3332 (
            .O(N__14734),
            .I(N__14710));
    LocalMux I__3331 (
            .O(N__14721),
            .I(N__14707));
    InMux I__3330 (
            .O(N__14720),
            .I(N__14702));
    InMux I__3329 (
            .O(N__14719),
            .I(N__14702));
    Span4Mux_v I__3328 (
            .O(N__14716),
            .I(N__14699));
    Span4Mux_s3_h I__3327 (
            .O(N__14713),
            .I(N__14696));
    LocalMux I__3326 (
            .O(N__14710),
            .I(N__14693));
    Span4Mux_v I__3325 (
            .O(N__14707),
            .I(N__14686));
    LocalMux I__3324 (
            .O(N__14702),
            .I(N__14686));
    Span4Mux_h I__3323 (
            .O(N__14699),
            .I(N__14686));
    Odrv4 I__3322 (
            .O(N__14696),
            .I(Lab_UT_di_Sones_2));
    Odrv12 I__3321 (
            .O(N__14693),
            .I(Lab_UT_di_Sones_2));
    Odrv4 I__3320 (
            .O(N__14686),
            .I(Lab_UT_di_Sones_2));
    CascadeMux I__3319 (
            .O(N__14679),
            .I(N__14676));
    InMux I__3318 (
            .O(N__14676),
            .I(N__14668));
    CascadeMux I__3317 (
            .O(N__14675),
            .I(N__14665));
    CascadeMux I__3316 (
            .O(N__14674),
            .I(N__14661));
    CascadeMux I__3315 (
            .O(N__14673),
            .I(N__14658));
    CascadeMux I__3314 (
            .O(N__14672),
            .I(N__14655));
    CascadeMux I__3313 (
            .O(N__14671),
            .I(N__14652));
    LocalMux I__3312 (
            .O(N__14668),
            .I(N__14647));
    InMux I__3311 (
            .O(N__14665),
            .I(N__14638));
    InMux I__3310 (
            .O(N__14664),
            .I(N__14638));
    InMux I__3309 (
            .O(N__14661),
            .I(N__14638));
    InMux I__3308 (
            .O(N__14658),
            .I(N__14638));
    InMux I__3307 (
            .O(N__14655),
            .I(N__14634));
    InMux I__3306 (
            .O(N__14652),
            .I(N__14629));
    InMux I__3305 (
            .O(N__14651),
            .I(N__14629));
    InMux I__3304 (
            .O(N__14650),
            .I(N__14626));
    Span4Mux_h I__3303 (
            .O(N__14647),
            .I(N__14623));
    LocalMux I__3302 (
            .O(N__14638),
            .I(N__14620));
    CascadeMux I__3301 (
            .O(N__14637),
            .I(N__14616));
    LocalMux I__3300 (
            .O(N__14634),
            .I(N__14613));
    LocalMux I__3299 (
            .O(N__14629),
            .I(N__14610));
    LocalMux I__3298 (
            .O(N__14626),
            .I(N__14605));
    Span4Mux_h I__3297 (
            .O(N__14623),
            .I(N__14605));
    Span4Mux_h I__3296 (
            .O(N__14620),
            .I(N__14602));
    InMux I__3295 (
            .O(N__14619),
            .I(N__14597));
    InMux I__3294 (
            .O(N__14616),
            .I(N__14597));
    Span4Mux_v I__3293 (
            .O(N__14613),
            .I(N__14592));
    Span4Mux_h I__3292 (
            .O(N__14610),
            .I(N__14592));
    Sp12to4 I__3291 (
            .O(N__14605),
            .I(N__14587));
    Sp12to4 I__3290 (
            .O(N__14602),
            .I(N__14587));
    LocalMux I__3289 (
            .O(N__14597),
            .I(Lab_UT_di_Sones_3));
    Odrv4 I__3288 (
            .O(N__14592),
            .I(Lab_UT_di_Sones_3));
    Odrv12 I__3287 (
            .O(N__14587),
            .I(Lab_UT_di_Sones_3));
    InMux I__3286 (
            .O(N__14580),
            .I(N__14577));
    LocalMux I__3285 (
            .O(N__14577),
            .I(\uu2.un1_segment3_m0 ));
    InMux I__3284 (
            .O(N__14574),
            .I(N__14569));
    CascadeMux I__3283 (
            .O(N__14573),
            .I(N__14565));
    InMux I__3282 (
            .O(N__14572),
            .I(N__14562));
    LocalMux I__3281 (
            .O(N__14569),
            .I(N__14559));
    InMux I__3280 (
            .O(N__14568),
            .I(N__14551));
    InMux I__3279 (
            .O(N__14565),
            .I(N__14548));
    LocalMux I__3278 (
            .O(N__14562),
            .I(N__14545));
    Span4Mux_v I__3277 (
            .O(N__14559),
            .I(N__14542));
    InMux I__3276 (
            .O(N__14558),
            .I(N__14537));
    InMux I__3275 (
            .O(N__14557),
            .I(N__14537));
    InMux I__3274 (
            .O(N__14556),
            .I(N__14530));
    InMux I__3273 (
            .O(N__14555),
            .I(N__14530));
    InMux I__3272 (
            .O(N__14554),
            .I(N__14530));
    LocalMux I__3271 (
            .O(N__14551),
            .I(N__14527));
    LocalMux I__3270 (
            .O(N__14548),
            .I(\uu2.w_addr_displaying_fastZ0Z_6 ));
    Odrv4 I__3269 (
            .O(N__14545),
            .I(\uu2.w_addr_displaying_fastZ0Z_6 ));
    Odrv4 I__3268 (
            .O(N__14542),
            .I(\uu2.w_addr_displaying_fastZ0Z_6 ));
    LocalMux I__3267 (
            .O(N__14537),
            .I(\uu2.w_addr_displaying_fastZ0Z_6 ));
    LocalMux I__3266 (
            .O(N__14530),
            .I(\uu2.w_addr_displaying_fastZ0Z_6 ));
    Odrv4 I__3265 (
            .O(N__14527),
            .I(\uu2.w_addr_displaying_fastZ0Z_6 ));
    CascadeMux I__3264 (
            .O(N__14514),
            .I(L3_segment1_3_cascade_));
    InMux I__3263 (
            .O(N__14511),
            .I(N__14507));
    InMux I__3262 (
            .O(N__14510),
            .I(N__14504));
    LocalMux I__3261 (
            .O(N__14507),
            .I(N__14497));
    LocalMux I__3260 (
            .O(N__14504),
            .I(N__14494));
    InMux I__3259 (
            .O(N__14503),
            .I(N__14491));
    InMux I__3258 (
            .O(N__14502),
            .I(N__14484));
    InMux I__3257 (
            .O(N__14501),
            .I(N__14484));
    InMux I__3256 (
            .O(N__14500),
            .I(N__14484));
    Span4Mux_h I__3255 (
            .O(N__14497),
            .I(N__14481));
    Odrv4 I__3254 (
            .O(N__14494),
            .I(\uu2.w_addr_displaying_fastZ0Z_5 ));
    LocalMux I__3253 (
            .O(N__14491),
            .I(\uu2.w_addr_displaying_fastZ0Z_5 ));
    LocalMux I__3252 (
            .O(N__14484),
            .I(\uu2.w_addr_displaying_fastZ0Z_5 ));
    Odrv4 I__3251 (
            .O(N__14481),
            .I(\uu2.w_addr_displaying_fastZ0Z_5 ));
    InMux I__3250 (
            .O(N__14472),
            .I(N__14469));
    LocalMux I__3249 (
            .O(N__14469),
            .I(N__14466));
    Odrv4 I__3248 (
            .O(N__14466),
            .I(\uu2.w_addr_displaying_fast_RNIQD7R4Z0Z_5 ));
    InMux I__3247 (
            .O(N__14463),
            .I(N__14458));
    InMux I__3246 (
            .O(N__14462),
            .I(N__14455));
    InMux I__3245 (
            .O(N__14461),
            .I(N__14450));
    LocalMux I__3244 (
            .O(N__14458),
            .I(N__14447));
    LocalMux I__3243 (
            .O(N__14455),
            .I(N__14444));
    InMux I__3242 (
            .O(N__14454),
            .I(N__14439));
    InMux I__3241 (
            .O(N__14453),
            .I(N__14439));
    LocalMux I__3240 (
            .O(N__14450),
            .I(N__14434));
    Span4Mux_h I__3239 (
            .O(N__14447),
            .I(N__14434));
    Odrv4 I__3238 (
            .O(N__14444),
            .I(\uu2.N_315_1 ));
    LocalMux I__3237 (
            .O(N__14439),
            .I(\uu2.N_315_1 ));
    Odrv4 I__3236 (
            .O(N__14434),
            .I(\uu2.N_315_1 ));
    InMux I__3235 (
            .O(N__14427),
            .I(N__14422));
    InMux I__3234 (
            .O(N__14426),
            .I(N__14417));
    InMux I__3233 (
            .O(N__14425),
            .I(N__14417));
    LocalMux I__3232 (
            .O(N__14422),
            .I(N__14410));
    LocalMux I__3231 (
            .O(N__14417),
            .I(N__14410));
    InMux I__3230 (
            .O(N__14416),
            .I(N__14405));
    InMux I__3229 (
            .O(N__14415),
            .I(N__14405));
    Odrv4 I__3228 (
            .O(N__14410),
            .I(\uu2.w_addr_displaying_4_rep2_RNI75VMZ0 ));
    LocalMux I__3227 (
            .O(N__14405),
            .I(\uu2.w_addr_displaying_4_rep2_RNI75VMZ0 ));
    InMux I__3226 (
            .O(N__14400),
            .I(N__14392));
    InMux I__3225 (
            .O(N__14399),
            .I(N__14392));
    InMux I__3224 (
            .O(N__14398),
            .I(N__14387));
    InMux I__3223 (
            .O(N__14397),
            .I(N__14387));
    LocalMux I__3222 (
            .O(N__14392),
            .I(N__14381));
    LocalMux I__3221 (
            .O(N__14387),
            .I(N__14378));
    InMux I__3220 (
            .O(N__14386),
            .I(N__14373));
    InMux I__3219 (
            .O(N__14385),
            .I(N__14373));
    CascadeMux I__3218 (
            .O(N__14384),
            .I(N__14370));
    Span4Mux_v I__3217 (
            .O(N__14381),
            .I(N__14366));
    Span4Mux_h I__3216 (
            .O(N__14378),
            .I(N__14363));
    LocalMux I__3215 (
            .O(N__14373),
            .I(N__14360));
    InMux I__3214 (
            .O(N__14370),
            .I(N__14355));
    InMux I__3213 (
            .O(N__14369),
            .I(N__14355));
    Odrv4 I__3212 (
            .O(N__14366),
            .I(\uu2.un1_segment3_m5 ));
    Odrv4 I__3211 (
            .O(N__14363),
            .I(\uu2.un1_segment3_m5 ));
    Odrv4 I__3210 (
            .O(N__14360),
            .I(\uu2.un1_segment3_m5 ));
    LocalMux I__3209 (
            .O(N__14355),
            .I(\uu2.un1_segment3_m5 ));
    InMux I__3208 (
            .O(N__14346),
            .I(N__14343));
    LocalMux I__3207 (
            .O(N__14343),
            .I(\uu2.N_813_0 ));
    InMux I__3206 (
            .O(N__14340),
            .I(N__14337));
    LocalMux I__3205 (
            .O(N__14337),
            .I(N__14334));
    Odrv12 I__3204 (
            .O(N__14334),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_59 ));
    CascadeMux I__3203 (
            .O(N__14331),
            .I(N__14328));
    InMux I__3202 (
            .O(N__14328),
            .I(N__14325));
    LocalMux I__3201 (
            .O(N__14325),
            .I(N__14322));
    Odrv12 I__3200 (
            .O(N__14322),
            .I(\uu2.segment2_m_2Z0Z_5 ));
    InMux I__3199 (
            .O(N__14319),
            .I(N__14316));
    LocalMux I__3198 (
            .O(N__14316),
            .I(\uu2.segment2_m_5 ));
    InMux I__3197 (
            .O(N__14313),
            .I(N__14309));
    InMux I__3196 (
            .O(N__14312),
            .I(N__14303));
    LocalMux I__3195 (
            .O(N__14309),
            .I(N__14300));
    InMux I__3194 (
            .O(N__14308),
            .I(N__14295));
    InMux I__3193 (
            .O(N__14307),
            .I(N__14295));
    InMux I__3192 (
            .O(N__14306),
            .I(N__14292));
    LocalMux I__3191 (
            .O(N__14303),
            .I(N__14289));
    Span4Mux_h I__3190 (
            .O(N__14300),
            .I(N__14279));
    LocalMux I__3189 (
            .O(N__14295),
            .I(N__14279));
    LocalMux I__3188 (
            .O(N__14292),
            .I(N__14274));
    Span4Mux_h I__3187 (
            .O(N__14289),
            .I(N__14274));
    InMux I__3186 (
            .O(N__14288),
            .I(N__14271));
    InMux I__3185 (
            .O(N__14287),
            .I(N__14262));
    InMux I__3184 (
            .O(N__14286),
            .I(N__14262));
    InMux I__3183 (
            .O(N__14285),
            .I(N__14262));
    InMux I__3182 (
            .O(N__14284),
            .I(N__14262));
    Odrv4 I__3181 (
            .O(N__14279),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    Odrv4 I__3180 (
            .O(N__14274),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__3179 (
            .O(N__14271),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__3178 (
            .O(N__14262),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    InMux I__3177 (
            .O(N__14253),
            .I(N__14250));
    LocalMux I__3176 (
            .O(N__14250),
            .I(N__14247));
    Span4Mux_v I__3175 (
            .O(N__14247),
            .I(N__14243));
    InMux I__3174 (
            .O(N__14246),
            .I(N__14240));
    Span4Mux_h I__3173 (
            .O(N__14243),
            .I(N__14235));
    LocalMux I__3172 (
            .O(N__14240),
            .I(N__14235));
    Span4Mux_v I__3171 (
            .O(N__14235),
            .I(N__14230));
    InMux I__3170 (
            .O(N__14234),
            .I(N__14227));
    InMux I__3169 (
            .O(N__14233),
            .I(N__14224));
    Span4Mux_h I__3168 (
            .O(N__14230),
            .I(N__14214));
    LocalMux I__3167 (
            .O(N__14227),
            .I(N__14214));
    LocalMux I__3166 (
            .O(N__14224),
            .I(N__14214));
    InMux I__3165 (
            .O(N__14223),
            .I(N__14209));
    InMux I__3164 (
            .O(N__14222),
            .I(N__14209));
    InMux I__3163 (
            .O(N__14221),
            .I(N__14206));
    Odrv4 I__3162 (
            .O(N__14214),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3161 (
            .O(N__14209),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3160 (
            .O(N__14206),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    InMux I__3159 (
            .O(N__14199),
            .I(N__14195));
    InMux I__3158 (
            .O(N__14198),
            .I(N__14192));
    LocalMux I__3157 (
            .O(N__14195),
            .I(N__14184));
    LocalMux I__3156 (
            .O(N__14192),
            .I(N__14181));
    InMux I__3155 (
            .O(N__14191),
            .I(N__14178));
    InMux I__3154 (
            .O(N__14190),
            .I(N__14171));
    InMux I__3153 (
            .O(N__14189),
            .I(N__14171));
    InMux I__3152 (
            .O(N__14188),
            .I(N__14171));
    InMux I__3151 (
            .O(N__14187),
            .I(N__14168));
    Span4Mux_v I__3150 (
            .O(N__14184),
            .I(N__14162));
    Span4Mux_v I__3149 (
            .O(N__14181),
            .I(N__14162));
    LocalMux I__3148 (
            .O(N__14178),
            .I(N__14155));
    LocalMux I__3147 (
            .O(N__14171),
            .I(N__14150));
    LocalMux I__3146 (
            .O(N__14168),
            .I(N__14150));
    InMux I__3145 (
            .O(N__14167),
            .I(N__14147));
    Span4Mux_h I__3144 (
            .O(N__14162),
            .I(N__14144));
    InMux I__3143 (
            .O(N__14161),
            .I(N__14135));
    InMux I__3142 (
            .O(N__14160),
            .I(N__14135));
    InMux I__3141 (
            .O(N__14159),
            .I(N__14135));
    InMux I__3140 (
            .O(N__14158),
            .I(N__14135));
    Span4Mux_h I__3139 (
            .O(N__14155),
            .I(N__14130));
    Span4Mux_v I__3138 (
            .O(N__14150),
            .I(N__14130));
    LocalMux I__3137 (
            .O(N__14147),
            .I(Lab_UT_di_Stens_2));
    Odrv4 I__3136 (
            .O(N__14144),
            .I(Lab_UT_di_Stens_2));
    LocalMux I__3135 (
            .O(N__14135),
            .I(Lab_UT_di_Stens_2));
    Odrv4 I__3134 (
            .O(N__14130),
            .I(Lab_UT_di_Stens_2));
    CascadeMux I__3133 (
            .O(N__14121),
            .I(N__14117));
    CascadeMux I__3132 (
            .O(N__14120),
            .I(N__14114));
    InMux I__3131 (
            .O(N__14117),
            .I(N__14107));
    InMux I__3130 (
            .O(N__14114),
            .I(N__14104));
    CascadeMux I__3129 (
            .O(N__14113),
            .I(N__14101));
    CascadeMux I__3128 (
            .O(N__14112),
            .I(N__14098));
    CascadeMux I__3127 (
            .O(N__14111),
            .I(N__14095));
    CascadeMux I__3126 (
            .O(N__14110),
            .I(N__14092));
    LocalMux I__3125 (
            .O(N__14107),
            .I(N__14083));
    LocalMux I__3124 (
            .O(N__14104),
            .I(N__14083));
    InMux I__3123 (
            .O(N__14101),
            .I(N__14080));
    InMux I__3122 (
            .O(N__14098),
            .I(N__14075));
    InMux I__3121 (
            .O(N__14095),
            .I(N__14075));
    InMux I__3120 (
            .O(N__14092),
            .I(N__14072));
    CascadeMux I__3119 (
            .O(N__14091),
            .I(N__14067));
    CascadeMux I__3118 (
            .O(N__14090),
            .I(N__14064));
    CascadeMux I__3117 (
            .O(N__14089),
            .I(N__14061));
    CascadeMux I__3116 (
            .O(N__14088),
            .I(N__14058));
    Span4Mux_v I__3115 (
            .O(N__14083),
            .I(N__14055));
    LocalMux I__3114 (
            .O(N__14080),
            .I(N__14048));
    LocalMux I__3113 (
            .O(N__14075),
            .I(N__14048));
    LocalMux I__3112 (
            .O(N__14072),
            .I(N__14048));
    InMux I__3111 (
            .O(N__14071),
            .I(N__14043));
    InMux I__3110 (
            .O(N__14070),
            .I(N__14043));
    InMux I__3109 (
            .O(N__14067),
            .I(N__14036));
    InMux I__3108 (
            .O(N__14064),
            .I(N__14036));
    InMux I__3107 (
            .O(N__14061),
            .I(N__14036));
    InMux I__3106 (
            .O(N__14058),
            .I(N__14033));
    Span4Mux_h I__3105 (
            .O(N__14055),
            .I(N__14028));
    Span4Mux_v I__3104 (
            .O(N__14048),
            .I(N__14028));
    LocalMux I__3103 (
            .O(N__14043),
            .I(Lab_UT_di_Stens_3));
    LocalMux I__3102 (
            .O(N__14036),
            .I(Lab_UT_di_Stens_3));
    LocalMux I__3101 (
            .O(N__14033),
            .I(Lab_UT_di_Stens_3));
    Odrv4 I__3100 (
            .O(N__14028),
            .I(Lab_UT_di_Stens_3));
    InMux I__3099 (
            .O(N__14019),
            .I(N__14016));
    LocalMux I__3098 (
            .O(N__14016),
            .I(\uu2.un1_segment3_m5_amZ0 ));
    InMux I__3097 (
            .O(N__14013),
            .I(N__14007));
    InMux I__3096 (
            .O(N__14012),
            .I(N__14004));
    InMux I__3095 (
            .O(N__14011),
            .I(N__14001));
    InMux I__3094 (
            .O(N__14010),
            .I(N__13998));
    LocalMux I__3093 (
            .O(N__14007),
            .I(N__13990));
    LocalMux I__3092 (
            .O(N__14004),
            .I(N__13990));
    LocalMux I__3091 (
            .O(N__14001),
            .I(N__13987));
    LocalMux I__3090 (
            .O(N__13998),
            .I(N__13984));
    InMux I__3089 (
            .O(N__13997),
            .I(N__13980));
    InMux I__3088 (
            .O(N__13996),
            .I(N__13977));
    InMux I__3087 (
            .O(N__13995),
            .I(N__13974));
    Span4Mux_v I__3086 (
            .O(N__13990),
            .I(N__13969));
    Span4Mux_v I__3085 (
            .O(N__13987),
            .I(N__13966));
    Span4Mux_h I__3084 (
            .O(N__13984),
            .I(N__13963));
    InMux I__3083 (
            .O(N__13983),
            .I(N__13960));
    LocalMux I__3082 (
            .O(N__13980),
            .I(N__13957));
    LocalMux I__3081 (
            .O(N__13977),
            .I(N__13952));
    LocalMux I__3080 (
            .O(N__13974),
            .I(N__13952));
    InMux I__3079 (
            .O(N__13973),
            .I(N__13949));
    InMux I__3078 (
            .O(N__13972),
            .I(N__13946));
    Odrv4 I__3077 (
            .O(N__13969),
            .I(\uu2.N_290_0_i_0 ));
    Odrv4 I__3076 (
            .O(N__13966),
            .I(\uu2.N_290_0_i_0 ));
    Odrv4 I__3075 (
            .O(N__13963),
            .I(\uu2.N_290_0_i_0 ));
    LocalMux I__3074 (
            .O(N__13960),
            .I(\uu2.N_290_0_i_0 ));
    Odrv4 I__3073 (
            .O(N__13957),
            .I(\uu2.N_290_0_i_0 ));
    Odrv4 I__3072 (
            .O(N__13952),
            .I(\uu2.N_290_0_i_0 ));
    LocalMux I__3071 (
            .O(N__13949),
            .I(\uu2.N_290_0_i_0 ));
    LocalMux I__3070 (
            .O(N__13946),
            .I(\uu2.N_290_0_i_0 ));
    CascadeMux I__3069 (
            .O(N__13929),
            .I(N__13926));
    InMux I__3068 (
            .O(N__13926),
            .I(N__13920));
    InMux I__3067 (
            .O(N__13925),
            .I(N__13920));
    LocalMux I__3066 (
            .O(N__13920),
            .I(N__13910));
    InMux I__3065 (
            .O(N__13919),
            .I(N__13903));
    InMux I__3064 (
            .O(N__13918),
            .I(N__13903));
    InMux I__3063 (
            .O(N__13917),
            .I(N__13903));
    CascadeMux I__3062 (
            .O(N__13916),
            .I(N__13900));
    InMux I__3061 (
            .O(N__13915),
            .I(N__13895));
    InMux I__3060 (
            .O(N__13914),
            .I(N__13895));
    CascadeMux I__3059 (
            .O(N__13913),
            .I(N__13892));
    Span4Mux_h I__3058 (
            .O(N__13910),
            .I(N__13889));
    LocalMux I__3057 (
            .O(N__13903),
            .I(N__13886));
    InMux I__3056 (
            .O(N__13900),
            .I(N__13883));
    LocalMux I__3055 (
            .O(N__13895),
            .I(N__13880));
    InMux I__3054 (
            .O(N__13892),
            .I(N__13877));
    Sp12to4 I__3053 (
            .O(N__13889),
            .I(N__13874));
    Span4Mux_v I__3052 (
            .O(N__13886),
            .I(N__13871));
    LocalMux I__3051 (
            .O(N__13883),
            .I(N__13866));
    Span4Mux_h I__3050 (
            .O(N__13880),
            .I(N__13866));
    LocalMux I__3049 (
            .O(N__13877),
            .I(\uu2.un436_ci ));
    Odrv12 I__3048 (
            .O(N__13874),
            .I(\uu2.un436_ci ));
    Odrv4 I__3047 (
            .O(N__13871),
            .I(\uu2.un436_ci ));
    Odrv4 I__3046 (
            .O(N__13866),
            .I(\uu2.un436_ci ));
    CascadeMux I__3045 (
            .O(N__13857),
            .I(N__13853));
    InMux I__3044 (
            .O(N__13856),
            .I(N__13848));
    InMux I__3043 (
            .O(N__13853),
            .I(N__13844));
    InMux I__3042 (
            .O(N__13852),
            .I(N__13838));
    InMux I__3041 (
            .O(N__13851),
            .I(N__13838));
    LocalMux I__3040 (
            .O(N__13848),
            .I(N__13835));
    InMux I__3039 (
            .O(N__13847),
            .I(N__13832));
    LocalMux I__3038 (
            .O(N__13844),
            .I(N__13829));
    CascadeMux I__3037 (
            .O(N__13843),
            .I(N__13823));
    LocalMux I__3036 (
            .O(N__13838),
            .I(N__13813));
    Span4Mux_v I__3035 (
            .O(N__13835),
            .I(N__13813));
    LocalMux I__3034 (
            .O(N__13832),
            .I(N__13813));
    Span4Mux_s3_h I__3033 (
            .O(N__13829),
            .I(N__13813));
    InMux I__3032 (
            .O(N__13828),
            .I(N__13808));
    InMux I__3031 (
            .O(N__13827),
            .I(N__13808));
    InMux I__3030 (
            .O(N__13826),
            .I(N__13805));
    InMux I__3029 (
            .O(N__13823),
            .I(N__13800));
    InMux I__3028 (
            .O(N__13822),
            .I(N__13800));
    Odrv4 I__3027 (
            .O(N__13813),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__3026 (
            .O(N__13808),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__3025 (
            .O(N__13805),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__3024 (
            .O(N__13800),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    InMux I__3023 (
            .O(N__13791),
            .I(N__13788));
    LocalMux I__3022 (
            .O(N__13788),
            .I(N__13785));
    Odrv12 I__3021 (
            .O(N__13785),
            .I(\uu2.un1_w_addr_displaying_35_0 ));
    InMux I__3020 (
            .O(N__13782),
            .I(N__13776));
    InMux I__3019 (
            .O(N__13781),
            .I(N__13772));
    CascadeMux I__3018 (
            .O(N__13780),
            .I(N__13766));
    InMux I__3017 (
            .O(N__13779),
            .I(N__13759));
    LocalMux I__3016 (
            .O(N__13776),
            .I(N__13753));
    InMux I__3015 (
            .O(N__13775),
            .I(N__13750));
    LocalMux I__3014 (
            .O(N__13772),
            .I(N__13747));
    InMux I__3013 (
            .O(N__13771),
            .I(N__13744));
    InMux I__3012 (
            .O(N__13770),
            .I(N__13737));
    InMux I__3011 (
            .O(N__13769),
            .I(N__13737));
    InMux I__3010 (
            .O(N__13766),
            .I(N__13737));
    InMux I__3009 (
            .O(N__13765),
            .I(N__13732));
    InMux I__3008 (
            .O(N__13764),
            .I(N__13732));
    InMux I__3007 (
            .O(N__13763),
            .I(N__13729));
    InMux I__3006 (
            .O(N__13762),
            .I(N__13726));
    LocalMux I__3005 (
            .O(N__13759),
            .I(N__13723));
    InMux I__3004 (
            .O(N__13758),
            .I(N__13718));
    InMux I__3003 (
            .O(N__13757),
            .I(N__13718));
    InMux I__3002 (
            .O(N__13756),
            .I(N__13715));
    Span4Mux_h I__3001 (
            .O(N__13753),
            .I(N__13708));
    LocalMux I__3000 (
            .O(N__13750),
            .I(N__13708));
    Span4Mux_h I__2999 (
            .O(N__13747),
            .I(N__13708));
    LocalMux I__2998 (
            .O(N__13744),
            .I(N__13705));
    LocalMux I__2997 (
            .O(N__13737),
            .I(N__13694));
    LocalMux I__2996 (
            .O(N__13732),
            .I(N__13694));
    LocalMux I__2995 (
            .O(N__13729),
            .I(N__13694));
    LocalMux I__2994 (
            .O(N__13726),
            .I(N__13694));
    Span4Mux_h I__2993 (
            .O(N__13723),
            .I(N__13694));
    LocalMux I__2992 (
            .O(N__13718),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2991 (
            .O(N__13715),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2990 (
            .O(N__13708),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2989 (
            .O(N__13705),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2988 (
            .O(N__13694),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    CascadeMux I__2987 (
            .O(N__13683),
            .I(\uu2.un1_w_addr_displaying_35_0_cascade_ ));
    InMux I__2986 (
            .O(N__13680),
            .I(N__13676));
    InMux I__2985 (
            .O(N__13679),
            .I(N__13673));
    LocalMux I__2984 (
            .O(N__13676),
            .I(\uu2.un1_w_addr_displaying_inv_2 ));
    LocalMux I__2983 (
            .O(N__13673),
            .I(\uu2.un1_w_addr_displaying_inv_2 ));
    CascadeMux I__2982 (
            .O(N__13668),
            .I(\uu2.N_813_0_cascade_ ));
    InMux I__2981 (
            .O(N__13665),
            .I(N__13662));
    LocalMux I__2980 (
            .O(N__13662),
            .I(N__13659));
    Odrv12 I__2979 (
            .O(N__13659),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_58 ));
    InMux I__2978 (
            .O(N__13656),
            .I(N__13649));
    InMux I__2977 (
            .O(N__13655),
            .I(N__13649));
    InMux I__2976 (
            .O(N__13654),
            .I(N__13646));
    LocalMux I__2975 (
            .O(N__13649),
            .I(N__13641));
    LocalMux I__2974 (
            .O(N__13646),
            .I(N__13641));
    Odrv12 I__2973 (
            .O(N__13641),
            .I(\Lab_UT.didpuu0.countEnMones ));
    InMux I__2972 (
            .O(N__13638),
            .I(N__13635));
    LocalMux I__2971 (
            .O(N__13635),
            .I(N__13632));
    Span4Mux_v I__2970 (
            .O(N__13632),
            .I(N__13629));
    Odrv4 I__2969 (
            .O(N__13629),
            .I(\uu2.un1_segment3_m5_bmZ0 ));
    InMux I__2968 (
            .O(N__13626),
            .I(N__13623));
    LocalMux I__2967 (
            .O(N__13623),
            .I(N__13619));
    InMux I__2966 (
            .O(N__13622),
            .I(N__13616));
    Span4Mux_v I__2965 (
            .O(N__13619),
            .I(N__13612));
    LocalMux I__2964 (
            .O(N__13616),
            .I(N__13609));
    InMux I__2963 (
            .O(N__13615),
            .I(N__13606));
    Odrv4 I__2962 (
            .O(N__13612),
            .I(bu_rx_data_1));
    Odrv12 I__2961 (
            .O(N__13609),
            .I(bu_rx_data_1));
    LocalMux I__2960 (
            .O(N__13606),
            .I(bu_rx_data_1));
    InMux I__2959 (
            .O(N__13599),
            .I(N__13596));
    LocalMux I__2958 (
            .O(N__13596),
            .I(N__13593));
    Sp12to4 I__2957 (
            .O(N__13593),
            .I(N__13589));
    InMux I__2956 (
            .O(N__13592),
            .I(N__13586));
    Span12Mux_s11_v I__2955 (
            .O(N__13589),
            .I(N__13581));
    LocalMux I__2954 (
            .O(N__13586),
            .I(N__13581));
    Odrv12 I__2953 (
            .O(N__13581),
            .I(bu_rx_data_0));
    CEMux I__2952 (
            .O(N__13578),
            .I(N__13574));
    CEMux I__2951 (
            .O(N__13577),
            .I(N__13571));
    LocalMux I__2950 (
            .O(N__13574),
            .I(N__13567));
    LocalMux I__2949 (
            .O(N__13571),
            .I(N__13564));
    CEMux I__2948 (
            .O(N__13570),
            .I(N__13561));
    Span4Mux_h I__2947 (
            .O(N__13567),
            .I(N__13554));
    Span4Mux_h I__2946 (
            .O(N__13564),
            .I(N__13554));
    LocalMux I__2945 (
            .O(N__13561),
            .I(N__13554));
    Span4Mux_h I__2944 (
            .O(N__13554),
            .I(N__13551));
    Odrv4 I__2943 (
            .O(N__13551),
            .I(\buart.Z_rx.N_41_i ));
    ClkMux I__2942 (
            .O(N__13548),
            .I(N__13350));
    ClkMux I__2941 (
            .O(N__13547),
            .I(N__13350));
    ClkMux I__2940 (
            .O(N__13546),
            .I(N__13350));
    ClkMux I__2939 (
            .O(N__13545),
            .I(N__13350));
    ClkMux I__2938 (
            .O(N__13544),
            .I(N__13350));
    ClkMux I__2937 (
            .O(N__13543),
            .I(N__13350));
    ClkMux I__2936 (
            .O(N__13542),
            .I(N__13350));
    ClkMux I__2935 (
            .O(N__13541),
            .I(N__13350));
    ClkMux I__2934 (
            .O(N__13540),
            .I(N__13350));
    ClkMux I__2933 (
            .O(N__13539),
            .I(N__13350));
    ClkMux I__2932 (
            .O(N__13538),
            .I(N__13350));
    ClkMux I__2931 (
            .O(N__13537),
            .I(N__13350));
    ClkMux I__2930 (
            .O(N__13536),
            .I(N__13350));
    ClkMux I__2929 (
            .O(N__13535),
            .I(N__13350));
    ClkMux I__2928 (
            .O(N__13534),
            .I(N__13350));
    ClkMux I__2927 (
            .O(N__13533),
            .I(N__13350));
    ClkMux I__2926 (
            .O(N__13532),
            .I(N__13350));
    ClkMux I__2925 (
            .O(N__13531),
            .I(N__13350));
    ClkMux I__2924 (
            .O(N__13530),
            .I(N__13350));
    ClkMux I__2923 (
            .O(N__13529),
            .I(N__13350));
    ClkMux I__2922 (
            .O(N__13528),
            .I(N__13350));
    ClkMux I__2921 (
            .O(N__13527),
            .I(N__13350));
    ClkMux I__2920 (
            .O(N__13526),
            .I(N__13350));
    ClkMux I__2919 (
            .O(N__13525),
            .I(N__13350));
    ClkMux I__2918 (
            .O(N__13524),
            .I(N__13350));
    ClkMux I__2917 (
            .O(N__13523),
            .I(N__13350));
    ClkMux I__2916 (
            .O(N__13522),
            .I(N__13350));
    ClkMux I__2915 (
            .O(N__13521),
            .I(N__13350));
    ClkMux I__2914 (
            .O(N__13520),
            .I(N__13350));
    ClkMux I__2913 (
            .O(N__13519),
            .I(N__13350));
    ClkMux I__2912 (
            .O(N__13518),
            .I(N__13350));
    ClkMux I__2911 (
            .O(N__13517),
            .I(N__13350));
    ClkMux I__2910 (
            .O(N__13516),
            .I(N__13350));
    ClkMux I__2909 (
            .O(N__13515),
            .I(N__13350));
    ClkMux I__2908 (
            .O(N__13514),
            .I(N__13350));
    ClkMux I__2907 (
            .O(N__13513),
            .I(N__13350));
    ClkMux I__2906 (
            .O(N__13512),
            .I(N__13350));
    ClkMux I__2905 (
            .O(N__13511),
            .I(N__13350));
    ClkMux I__2904 (
            .O(N__13510),
            .I(N__13350));
    ClkMux I__2903 (
            .O(N__13509),
            .I(N__13350));
    ClkMux I__2902 (
            .O(N__13508),
            .I(N__13350));
    ClkMux I__2901 (
            .O(N__13507),
            .I(N__13350));
    ClkMux I__2900 (
            .O(N__13506),
            .I(N__13350));
    ClkMux I__2899 (
            .O(N__13505),
            .I(N__13350));
    ClkMux I__2898 (
            .O(N__13504),
            .I(N__13350));
    ClkMux I__2897 (
            .O(N__13503),
            .I(N__13350));
    ClkMux I__2896 (
            .O(N__13502),
            .I(N__13350));
    ClkMux I__2895 (
            .O(N__13501),
            .I(N__13350));
    ClkMux I__2894 (
            .O(N__13500),
            .I(N__13350));
    ClkMux I__2893 (
            .O(N__13499),
            .I(N__13350));
    ClkMux I__2892 (
            .O(N__13498),
            .I(N__13350));
    ClkMux I__2891 (
            .O(N__13497),
            .I(N__13350));
    ClkMux I__2890 (
            .O(N__13496),
            .I(N__13350));
    ClkMux I__2889 (
            .O(N__13495),
            .I(N__13350));
    ClkMux I__2888 (
            .O(N__13494),
            .I(N__13350));
    ClkMux I__2887 (
            .O(N__13493),
            .I(N__13350));
    ClkMux I__2886 (
            .O(N__13492),
            .I(N__13350));
    ClkMux I__2885 (
            .O(N__13491),
            .I(N__13350));
    ClkMux I__2884 (
            .O(N__13490),
            .I(N__13350));
    ClkMux I__2883 (
            .O(N__13489),
            .I(N__13350));
    ClkMux I__2882 (
            .O(N__13488),
            .I(N__13350));
    ClkMux I__2881 (
            .O(N__13487),
            .I(N__13350));
    ClkMux I__2880 (
            .O(N__13486),
            .I(N__13350));
    ClkMux I__2879 (
            .O(N__13485),
            .I(N__13350));
    ClkMux I__2878 (
            .O(N__13484),
            .I(N__13350));
    ClkMux I__2877 (
            .O(N__13483),
            .I(N__13350));
    GlobalMux I__2876 (
            .O(N__13350),
            .I(N__13347));
    gio2CtrlBuf I__2875 (
            .O(N__13347),
            .I(clk_g));
    CascadeMux I__2874 (
            .O(N__13344),
            .I(N__13341));
    InMux I__2873 (
            .O(N__13341),
            .I(N__13338));
    LocalMux I__2872 (
            .O(N__13338),
            .I(N__13335));
    Span12Mux_s4_h I__2871 (
            .O(N__13335),
            .I(N__13331));
    InMux I__2870 (
            .O(N__13334),
            .I(N__13328));
    Odrv12 I__2869 (
            .O(N__13331),
            .I(\Lab_UT.sec_clkD ));
    LocalMux I__2868 (
            .O(N__13328),
            .I(\Lab_UT.sec_clkD ));
    InMux I__2867 (
            .O(N__13323),
            .I(N__13318));
    InMux I__2866 (
            .O(N__13322),
            .I(N__13313));
    InMux I__2865 (
            .O(N__13321),
            .I(N__13313));
    LocalMux I__2864 (
            .O(N__13318),
            .I(N__13308));
    LocalMux I__2863 (
            .O(N__13313),
            .I(N__13308));
    Span4Mux_v I__2862 (
            .O(N__13308),
            .I(N__13303));
    InMux I__2861 (
            .O(N__13307),
            .I(N__13298));
    InMux I__2860 (
            .O(N__13306),
            .I(N__13298));
    Odrv4 I__2859 (
            .O(N__13303),
            .I(\Lab_UT.didpuu0.clkSecStrbZ0 ));
    LocalMux I__2858 (
            .O(N__13298),
            .I(\Lab_UT.didpuu0.clkSecStrbZ0 ));
    InMux I__2857 (
            .O(N__13293),
            .I(N__13290));
    LocalMux I__2856 (
            .O(N__13290),
            .I(N__13287));
    Span4Mux_h I__2855 (
            .O(N__13287),
            .I(N__13284));
    Odrv4 I__2854 (
            .O(N__13284),
            .I(L3_segment3_2));
    CascadeMux I__2853 (
            .O(N__13281),
            .I(L3_segment2_4_cascade_));
    InMux I__2852 (
            .O(N__13278),
            .I(N__13275));
    LocalMux I__2851 (
            .O(N__13275),
            .I(N__13272));
    Span4Mux_h I__2850 (
            .O(N__13272),
            .I(N__13269));
    Odrv4 I__2849 (
            .O(N__13269),
            .I(\uu2.segment2_m_1Z0Z_6 ));
    CascadeMux I__2848 (
            .O(N__13266),
            .I(\Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMUZ0Z_0_cascade_ ));
    IoInMux I__2847 (
            .O(N__13263),
            .I(N__13260));
    LocalMux I__2846 (
            .O(N__13260),
            .I(N__13257));
    Span4Mux_s3_h I__2845 (
            .O(N__13257),
            .I(N__13254));
    Odrv4 I__2844 (
            .O(N__13254),
            .I(led_c_3));
    InMux I__2843 (
            .O(N__13251),
            .I(N__13248));
    LocalMux I__2842 (
            .O(N__13248),
            .I(\Lab_UT.didpuu0.ledDisp00.selLed_RNI67CIZ0Z_0 ));
    CascadeMux I__2841 (
            .O(N__13245),
            .I(N__13241));
    CascadeMux I__2840 (
            .O(N__13244),
            .I(N__13238));
    InMux I__2839 (
            .O(N__13241),
            .I(N__13233));
    InMux I__2838 (
            .O(N__13238),
            .I(N__13233));
    LocalMux I__2837 (
            .O(N__13233),
            .I(N__13230));
    Span4Mux_v I__2836 (
            .O(N__13230),
            .I(N__13226));
    InMux I__2835 (
            .O(N__13229),
            .I(N__13223));
    Odrv4 I__2834 (
            .O(N__13226),
            .I(\Lab_UT.un11_segmentUQ_1 ));
    LocalMux I__2833 (
            .O(N__13223),
            .I(\Lab_UT.un11_segmentUQ_1 ));
    CascadeMux I__2832 (
            .O(N__13218),
            .I(\Lab_UT.didpuu0.countEnMtens_0_a4_0_cascade_ ));
    InMux I__2831 (
            .O(N__13215),
            .I(N__13211));
    InMux I__2830 (
            .O(N__13214),
            .I(N__13208));
    LocalMux I__2829 (
            .O(N__13211),
            .I(N__13205));
    LocalMux I__2828 (
            .O(N__13208),
            .I(N__13202));
    Span4Mux_v I__2827 (
            .O(N__13205),
            .I(N__13199));
    Span4Mux_v I__2826 (
            .O(N__13202),
            .I(N__13194));
    Span4Mux_h I__2825 (
            .O(N__13199),
            .I(N__13194));
    Odrv4 I__2824 (
            .O(N__13194),
            .I(\Lab_UT.didpuu0.countEnMtens_0_a4_1 ));
    CascadeMux I__2823 (
            .O(N__13191),
            .I(\Lab_UT.didpuu0.countEnMtens_0_a4_1_cascade_ ));
    InMux I__2822 (
            .O(N__13188),
            .I(N__13185));
    LocalMux I__2821 (
            .O(N__13185),
            .I(N__13180));
    InMux I__2820 (
            .O(N__13184),
            .I(N__13174));
    InMux I__2819 (
            .O(N__13183),
            .I(N__13171));
    Span4Mux_v I__2818 (
            .O(N__13180),
            .I(N__13168));
    InMux I__2817 (
            .O(N__13179),
            .I(N__13161));
    InMux I__2816 (
            .O(N__13178),
            .I(N__13161));
    InMux I__2815 (
            .O(N__13177),
            .I(N__13161));
    LocalMux I__2814 (
            .O(N__13174),
            .I(\Lab_UT.didpuu0.countEnStens ));
    LocalMux I__2813 (
            .O(N__13171),
            .I(\Lab_UT.didpuu0.countEnStens ));
    Odrv4 I__2812 (
            .O(N__13168),
            .I(\Lab_UT.didpuu0.countEnStens ));
    LocalMux I__2811 (
            .O(N__13161),
            .I(\Lab_UT.didpuu0.countEnStens ));
    InMux I__2810 (
            .O(N__13152),
            .I(N__13148));
    InMux I__2809 (
            .O(N__13151),
            .I(N__13145));
    LocalMux I__2808 (
            .O(N__13148),
            .I(N__13142));
    LocalMux I__2807 (
            .O(N__13145),
            .I(N__13139));
    Span4Mux_h I__2806 (
            .O(N__13142),
            .I(N__13136));
    Sp12to4 I__2805 (
            .O(N__13139),
            .I(N__13133));
    Span4Mux_v I__2804 (
            .O(N__13136),
            .I(N__13130));
    Odrv12 I__2803 (
            .O(N__13133),
            .I(\Lab_UT.didpuu0.countEnMtens ));
    Odrv4 I__2802 (
            .O(N__13130),
            .I(\Lab_UT.didpuu0.countEnMtens ));
    InMux I__2801 (
            .O(N__13125),
            .I(N__13122));
    LocalMux I__2800 (
            .O(N__13122),
            .I(\Lab_UT.un152_segmentUQ_1 ));
    CEMux I__2799 (
            .O(N__13119),
            .I(N__13116));
    LocalMux I__2798 (
            .O(N__13116),
            .I(N__13113));
    Span4Mux_v I__2797 (
            .O(N__13113),
            .I(N__13110));
    Odrv4 I__2796 (
            .O(N__13110),
            .I(\Lab_UT.didpuu0.didpstens.countEnStens_0 ));
    InMux I__2795 (
            .O(N__13107),
            .I(N__13104));
    LocalMux I__2794 (
            .O(N__13104),
            .I(\uu2.un1_segment4_3_bmZ0 ));
    CascadeMux I__2793 (
            .O(N__13101),
            .I(\uu2.un1_segment4_3_amZ0_cascade_ ));
    InMux I__2792 (
            .O(N__13098),
            .I(N__13095));
    LocalMux I__2791 (
            .O(N__13095),
            .I(\uu2.un1_segment4_9_ns_1 ));
    CascadeMux I__2790 (
            .O(N__13092),
            .I(\uu2.N_289_cascade_ ));
    InMux I__2789 (
            .O(N__13089),
            .I(N__13086));
    LocalMux I__2788 (
            .O(N__13086),
            .I(\uu2.w_addr_displaying_fast_RNIFU9M8Z0Z_8 ));
    InMux I__2787 (
            .O(N__13083),
            .I(N__13078));
    CascadeMux I__2786 (
            .O(N__13082),
            .I(N__13074));
    InMux I__2785 (
            .O(N__13081),
            .I(N__13071));
    LocalMux I__2784 (
            .O(N__13078),
            .I(N__13066));
    InMux I__2783 (
            .O(N__13077),
            .I(N__13061));
    InMux I__2782 (
            .O(N__13074),
            .I(N__13061));
    LocalMux I__2781 (
            .O(N__13071),
            .I(N__13057));
    InMux I__2780 (
            .O(N__13070),
            .I(N__13052));
    InMux I__2779 (
            .O(N__13069),
            .I(N__13052));
    Span4Mux_h I__2778 (
            .O(N__13066),
            .I(N__13047));
    LocalMux I__2777 (
            .O(N__13061),
            .I(N__13047));
    InMux I__2776 (
            .O(N__13060),
            .I(N__13044));
    Odrv4 I__2775 (
            .O(N__13057),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__2774 (
            .O(N__13052),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    Odrv4 I__2773 (
            .O(N__13047),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__2772 (
            .O(N__13044),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    CascadeMux I__2771 (
            .O(N__13035),
            .I(N__13032));
    InMux I__2770 (
            .O(N__13032),
            .I(N__13029));
    LocalMux I__2769 (
            .O(N__13029),
            .I(N__13026));
    Span4Mux_h I__2768 (
            .O(N__13026),
            .I(N__13023));
    Odrv4 I__2767 (
            .O(N__13023),
            .I(\uu2.N_1 ));
    InMux I__2766 (
            .O(N__13020),
            .I(N__13017));
    LocalMux I__2765 (
            .O(N__13017),
            .I(\uu2.w_addr_displaying_4_rep1_RNIAVDBZ0Z_0 ));
    InMux I__2764 (
            .O(N__13014),
            .I(N__13011));
    LocalMux I__2763 (
            .O(N__13011),
            .I(N__13008));
    Span4Mux_h I__2762 (
            .O(N__13008),
            .I(N__13005));
    Odrv4 I__2761 (
            .O(N__13005),
            .I(\uu2.w_addr_displaying_fast_RNIKFIEZ0Z_6 ));
    InMux I__2760 (
            .O(N__13002),
            .I(N__12999));
    LocalMux I__2759 (
            .O(N__12999),
            .I(N__12996));
    Span4Mux_h I__2758 (
            .O(N__12996),
            .I(N__12993));
    Odrv4 I__2757 (
            .O(N__12993),
            .I(\uu2.w_addr_displaying_fast_RNIN0TSZ0Z_4 ));
    InMux I__2756 (
            .O(N__12990),
            .I(N__12980));
    InMux I__2755 (
            .O(N__12989),
            .I(N__12980));
    InMux I__2754 (
            .O(N__12988),
            .I(N__12977));
    InMux I__2753 (
            .O(N__12987),
            .I(N__12970));
    InMux I__2752 (
            .O(N__12986),
            .I(N__12970));
    InMux I__2751 (
            .O(N__12985),
            .I(N__12970));
    LocalMux I__2750 (
            .O(N__12980),
            .I(\uu2.w_addr_displaying_fastZ0Z_4 ));
    LocalMux I__2749 (
            .O(N__12977),
            .I(\uu2.w_addr_displaying_fastZ0Z_4 ));
    LocalMux I__2748 (
            .O(N__12970),
            .I(\uu2.w_addr_displaying_fastZ0Z_4 ));
    CascadeMux I__2747 (
            .O(N__12963),
            .I(N__12958));
    InMux I__2746 (
            .O(N__12962),
            .I(N__12955));
    InMux I__2745 (
            .O(N__12961),
            .I(N__12949));
    InMux I__2744 (
            .O(N__12958),
            .I(N__12946));
    LocalMux I__2743 (
            .O(N__12955),
            .I(N__12943));
    InMux I__2742 (
            .O(N__12954),
            .I(N__12940));
    InMux I__2741 (
            .O(N__12953),
            .I(N__12935));
    InMux I__2740 (
            .O(N__12952),
            .I(N__12935));
    LocalMux I__2739 (
            .O(N__12949),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    LocalMux I__2738 (
            .O(N__12946),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    Odrv4 I__2737 (
            .O(N__12943),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    LocalMux I__2736 (
            .O(N__12940),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    LocalMux I__2735 (
            .O(N__12935),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    InMux I__2734 (
            .O(N__12924),
            .I(N__12921));
    LocalMux I__2733 (
            .O(N__12921),
            .I(\uu2.N_10_0 ));
    CascadeMux I__2732 (
            .O(N__12918),
            .I(N__12914));
    InMux I__2731 (
            .O(N__12917),
            .I(N__12911));
    InMux I__2730 (
            .O(N__12914),
            .I(N__12908));
    LocalMux I__2729 (
            .O(N__12911),
            .I(N__12905));
    LocalMux I__2728 (
            .O(N__12908),
            .I(N__12902));
    Span4Mux_h I__2727 (
            .O(N__12905),
            .I(N__12899));
    Span4Mux_h I__2726 (
            .O(N__12902),
            .I(N__12894));
    Span4Mux_v I__2725 (
            .O(N__12899),
            .I(N__12894));
    Odrv4 I__2724 (
            .O(N__12894),
            .I(\Lab_UT.didpuu0.didpsones.N_38 ));
    CascadeMux I__2723 (
            .O(N__12891),
            .I(N__12888));
    InMux I__2722 (
            .O(N__12888),
            .I(N__12885));
    LocalMux I__2721 (
            .O(N__12885),
            .I(N__12882));
    Span4Mux_v I__2720 (
            .O(N__12882),
            .I(N__12879));
    Span4Mux_s3_h I__2719 (
            .O(N__12879),
            .I(N__12876));
    Odrv4 I__2718 (
            .O(N__12876),
            .I(\Lab_UT.didpuu0.didpsones.N_32 ));
    InMux I__2717 (
            .O(N__12873),
            .I(N__12869));
    InMux I__2716 (
            .O(N__12872),
            .I(N__12865));
    LocalMux I__2715 (
            .O(N__12869),
            .I(N__12862));
    InMux I__2714 (
            .O(N__12868),
            .I(N__12859));
    LocalMux I__2713 (
            .O(N__12865),
            .I(N__12856));
    Span4Mux_h I__2712 (
            .O(N__12862),
            .I(N__12849));
    LocalMux I__2711 (
            .O(N__12859),
            .I(N__12849));
    Span4Mux_h I__2710 (
            .O(N__12856),
            .I(N__12849));
    Odrv4 I__2709 (
            .O(N__12849),
            .I(Lab_UT_dec0_un137_segmentUQ));
    CascadeMux I__2708 (
            .O(N__12846),
            .I(\uu2.segment1_m_2Z0Z_0_cascade_ ));
    CascadeMux I__2707 (
            .O(N__12843),
            .I(\uu2.segment1_m_0_cascade_ ));
    InMux I__2706 (
            .O(N__12840),
            .I(N__12831));
    InMux I__2705 (
            .O(N__12839),
            .I(N__12826));
    InMux I__2704 (
            .O(N__12838),
            .I(N__12826));
    InMux I__2703 (
            .O(N__12837),
            .I(N__12823));
    InMux I__2702 (
            .O(N__12836),
            .I(N__12820));
    InMux I__2701 (
            .O(N__12835),
            .I(N__12814));
    InMux I__2700 (
            .O(N__12834),
            .I(N__12814));
    LocalMux I__2699 (
            .O(N__12831),
            .I(N__12805));
    LocalMux I__2698 (
            .O(N__12826),
            .I(N__12805));
    LocalMux I__2697 (
            .O(N__12823),
            .I(N__12800));
    LocalMux I__2696 (
            .O(N__12820),
            .I(N__12800));
    InMux I__2695 (
            .O(N__12819),
            .I(N__12791));
    LocalMux I__2694 (
            .O(N__12814),
            .I(N__12788));
    InMux I__2693 (
            .O(N__12813),
            .I(N__12779));
    InMux I__2692 (
            .O(N__12812),
            .I(N__12779));
    InMux I__2691 (
            .O(N__12811),
            .I(N__12779));
    InMux I__2690 (
            .O(N__12810),
            .I(N__12779));
    Span4Mux_v I__2689 (
            .O(N__12805),
            .I(N__12774));
    Span4Mux_h I__2688 (
            .O(N__12800),
            .I(N__12774));
    InMux I__2687 (
            .O(N__12799),
            .I(N__12767));
    InMux I__2686 (
            .O(N__12798),
            .I(N__12767));
    InMux I__2685 (
            .O(N__12797),
            .I(N__12767));
    InMux I__2684 (
            .O(N__12796),
            .I(N__12764));
    InMux I__2683 (
            .O(N__12795),
            .I(N__12761));
    InMux I__2682 (
            .O(N__12794),
            .I(N__12758));
    LocalMux I__2681 (
            .O(N__12791),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2680 (
            .O(N__12788),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2679 (
            .O(N__12779),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2678 (
            .O(N__12774),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2677 (
            .O(N__12767),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2676 (
            .O(N__12764),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2675 (
            .O(N__12761),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2674 (
            .O(N__12758),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    InMux I__2673 (
            .O(N__12741),
            .I(N__12738));
    LocalMux I__2672 (
            .O(N__12738),
            .I(\uu2.segment3_m_6 ));
    CascadeMux I__2671 (
            .O(N__12735),
            .I(\uu2.un1_segment1_iv_0_cascade_ ));
    InMux I__2670 (
            .O(N__12732),
            .I(N__12724));
    InMux I__2669 (
            .O(N__12731),
            .I(N__12719));
    InMux I__2668 (
            .O(N__12730),
            .I(N__12719));
    CascadeMux I__2667 (
            .O(N__12729),
            .I(N__12716));
    CascadeMux I__2666 (
            .O(N__12728),
            .I(N__12712));
    CascadeMux I__2665 (
            .O(N__12727),
            .I(N__12709));
    LocalMux I__2664 (
            .O(N__12724),
            .I(N__12704));
    LocalMux I__2663 (
            .O(N__12719),
            .I(N__12704));
    InMux I__2662 (
            .O(N__12716),
            .I(N__12699));
    InMux I__2661 (
            .O(N__12715),
            .I(N__12699));
    InMux I__2660 (
            .O(N__12712),
            .I(N__12694));
    InMux I__2659 (
            .O(N__12709),
            .I(N__12694));
    Span4Mux_h I__2658 (
            .O(N__12704),
            .I(N__12691));
    LocalMux I__2657 (
            .O(N__12699),
            .I(N__12686));
    LocalMux I__2656 (
            .O(N__12694),
            .I(N__12686));
    Odrv4 I__2655 (
            .O(N__12691),
            .I(\uu2.un1_segment1_0 ));
    Odrv4 I__2654 (
            .O(N__12686),
            .I(\uu2.un1_segment1_0 ));
    InMux I__2653 (
            .O(N__12681),
            .I(N__12678));
    LocalMux I__2652 (
            .O(N__12678),
            .I(\uu2.un1_segment4_sn_N_61 ));
    CascadeMux I__2651 (
            .O(N__12675),
            .I(\uu2.w_addr_displaying_fast_RNI6N2KZ0Z_5_cascade_ ));
    InMux I__2650 (
            .O(N__12672),
            .I(N__12669));
    LocalMux I__2649 (
            .O(N__12669),
            .I(\uu2.w_addr_displaying_fast_RNID5QHZ0Z_5 ));
    InMux I__2648 (
            .O(N__12666),
            .I(N__12663));
    LocalMux I__2647 (
            .O(N__12663),
            .I(N__12660));
    Odrv4 I__2646 (
            .O(N__12660),
            .I(\uu2.un1_segment4_sn_N_39_0 ));
    InMux I__2645 (
            .O(N__12657),
            .I(N__12654));
    LocalMux I__2644 (
            .O(N__12654),
            .I(N__12651));
    Odrv12 I__2643 (
            .O(N__12651),
            .I(\uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4 ));
    CascadeMux I__2642 (
            .O(N__12648),
            .I(\uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4_cascade_ ));
    CascadeMux I__2641 (
            .O(N__12645),
            .I(N__12640));
    InMux I__2640 (
            .O(N__12644),
            .I(N__12635));
    InMux I__2639 (
            .O(N__12643),
            .I(N__12635));
    InMux I__2638 (
            .O(N__12640),
            .I(N__12632));
    LocalMux I__2637 (
            .O(N__12635),
            .I(N__12627));
    LocalMux I__2636 (
            .O(N__12632),
            .I(N__12624));
    InMux I__2635 (
            .O(N__12631),
            .I(N__12619));
    InMux I__2634 (
            .O(N__12630),
            .I(N__12619));
    Span4Mux_h I__2633 (
            .O(N__12627),
            .I(N__12614));
    Span4Mux_h I__2632 (
            .O(N__12624),
            .I(N__12609));
    LocalMux I__2631 (
            .O(N__12619),
            .I(N__12609));
    InMux I__2630 (
            .O(N__12618),
            .I(N__12604));
    InMux I__2629 (
            .O(N__12617),
            .I(N__12604));
    Odrv4 I__2628 (
            .O(N__12614),
            .I(\uu2.w_addr_displaying_RNILB202Z0Z_4 ));
    Odrv4 I__2627 (
            .O(N__12609),
            .I(\uu2.w_addr_displaying_RNILB202Z0Z_4 ));
    LocalMux I__2626 (
            .O(N__12604),
            .I(\uu2.w_addr_displaying_RNILB202Z0Z_4 ));
    InMux I__2625 (
            .O(N__12597),
            .I(N__12594));
    LocalMux I__2624 (
            .O(N__12594),
            .I(N__12591));
    Span4Mux_h I__2623 (
            .O(N__12591),
            .I(N__12588));
    Odrv4 I__2622 (
            .O(N__12588),
            .I(\uu2.N_92 ));
    CascadeMux I__2621 (
            .O(N__12585),
            .I(N__12582));
    InMux I__2620 (
            .O(N__12582),
            .I(N__12579));
    LocalMux I__2619 (
            .O(N__12579),
            .I(\uu2.w_addr_displaying_4_0_i_fast_6 ));
    InMux I__2618 (
            .O(N__12576),
            .I(N__12572));
    CascadeMux I__2617 (
            .O(N__12575),
            .I(N__12566));
    LocalMux I__2616 (
            .O(N__12572),
            .I(N__12558));
    InMux I__2615 (
            .O(N__12571),
            .I(N__12551));
    InMux I__2614 (
            .O(N__12570),
            .I(N__12551));
    InMux I__2613 (
            .O(N__12569),
            .I(N__12551));
    InMux I__2612 (
            .O(N__12566),
            .I(N__12548));
    InMux I__2611 (
            .O(N__12565),
            .I(N__12545));
    InMux I__2610 (
            .O(N__12564),
            .I(N__12540));
    InMux I__2609 (
            .O(N__12563),
            .I(N__12540));
    InMux I__2608 (
            .O(N__12562),
            .I(N__12535));
    InMux I__2607 (
            .O(N__12561),
            .I(N__12535));
    Span4Mux_h I__2606 (
            .O(N__12558),
            .I(N__12531));
    LocalMux I__2605 (
            .O(N__12551),
            .I(N__12528));
    LocalMux I__2604 (
            .O(N__12548),
            .I(N__12525));
    LocalMux I__2603 (
            .O(N__12545),
            .I(N__12516));
    LocalMux I__2602 (
            .O(N__12540),
            .I(N__12516));
    LocalMux I__2601 (
            .O(N__12535),
            .I(N__12516));
    InMux I__2600 (
            .O(N__12534),
            .I(N__12513));
    Span4Mux_h I__2599 (
            .O(N__12531),
            .I(N__12510));
    Span4Mux_v I__2598 (
            .O(N__12528),
            .I(N__12505));
    Span4Mux_h I__2597 (
            .O(N__12525),
            .I(N__12505));
    InMux I__2596 (
            .O(N__12524),
            .I(N__12500));
    InMux I__2595 (
            .O(N__12523),
            .I(N__12500));
    Span4Mux_v I__2594 (
            .O(N__12516),
            .I(N__12497));
    LocalMux I__2593 (
            .O(N__12513),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2592 (
            .O(N__12510),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2591 (
            .O(N__12505),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2590 (
            .O(N__12500),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2589 (
            .O(N__12497),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    CascadeMux I__2588 (
            .O(N__12486),
            .I(\uu2.un15_w_data_displaying_cascade_ ));
    CascadeMux I__2587 (
            .O(N__12483),
            .I(N__12479));
    CascadeMux I__2586 (
            .O(N__12482),
            .I(N__12472));
    InMux I__2585 (
            .O(N__12479),
            .I(N__12463));
    InMux I__2584 (
            .O(N__12478),
            .I(N__12451));
    InMux I__2583 (
            .O(N__12477),
            .I(N__12451));
    InMux I__2582 (
            .O(N__12476),
            .I(N__12451));
    InMux I__2581 (
            .O(N__12475),
            .I(N__12451));
    InMux I__2580 (
            .O(N__12472),
            .I(N__12448));
    InMux I__2579 (
            .O(N__12471),
            .I(N__12445));
    InMux I__2578 (
            .O(N__12470),
            .I(N__12440));
    InMux I__2577 (
            .O(N__12469),
            .I(N__12440));
    InMux I__2576 (
            .O(N__12468),
            .I(N__12433));
    InMux I__2575 (
            .O(N__12467),
            .I(N__12433));
    InMux I__2574 (
            .O(N__12466),
            .I(N__12433));
    LocalMux I__2573 (
            .O(N__12463),
            .I(N__12430));
    CascadeMux I__2572 (
            .O(N__12462),
            .I(N__12421));
    InMux I__2571 (
            .O(N__12461),
            .I(N__12415));
    InMux I__2570 (
            .O(N__12460),
            .I(N__12415));
    LocalMux I__2569 (
            .O(N__12451),
            .I(N__12412));
    LocalMux I__2568 (
            .O(N__12448),
            .I(N__12405));
    LocalMux I__2567 (
            .O(N__12445),
            .I(N__12405));
    LocalMux I__2566 (
            .O(N__12440),
            .I(N__12405));
    LocalMux I__2565 (
            .O(N__12433),
            .I(N__12400));
    Span4Mux_v I__2564 (
            .O(N__12430),
            .I(N__12400));
    InMux I__2563 (
            .O(N__12429),
            .I(N__12392));
    InMux I__2562 (
            .O(N__12428),
            .I(N__12392));
    InMux I__2561 (
            .O(N__12427),
            .I(N__12392));
    InMux I__2560 (
            .O(N__12426),
            .I(N__12389));
    InMux I__2559 (
            .O(N__12425),
            .I(N__12386));
    InMux I__2558 (
            .O(N__12424),
            .I(N__12379));
    InMux I__2557 (
            .O(N__12421),
            .I(N__12379));
    InMux I__2556 (
            .O(N__12420),
            .I(N__12379));
    LocalMux I__2555 (
            .O(N__12415),
            .I(N__12376));
    Span4Mux_v I__2554 (
            .O(N__12412),
            .I(N__12371));
    Span4Mux_v I__2553 (
            .O(N__12405),
            .I(N__12371));
    Span4Mux_h I__2552 (
            .O(N__12400),
            .I(N__12368));
    InMux I__2551 (
            .O(N__12399),
            .I(N__12365));
    LocalMux I__2550 (
            .O(N__12392),
            .I(N__12360));
    LocalMux I__2549 (
            .O(N__12389),
            .I(N__12360));
    LocalMux I__2548 (
            .O(N__12386),
            .I(\uu2.un19_w_addr_userZ0Z_0 ));
    LocalMux I__2547 (
            .O(N__12379),
            .I(\uu2.un19_w_addr_userZ0Z_0 ));
    Odrv4 I__2546 (
            .O(N__12376),
            .I(\uu2.un19_w_addr_userZ0Z_0 ));
    Odrv4 I__2545 (
            .O(N__12371),
            .I(\uu2.un19_w_addr_userZ0Z_0 ));
    Odrv4 I__2544 (
            .O(N__12368),
            .I(\uu2.un19_w_addr_userZ0Z_0 ));
    LocalMux I__2543 (
            .O(N__12365),
            .I(\uu2.un19_w_addr_userZ0Z_0 ));
    Odrv12 I__2542 (
            .O(N__12360),
            .I(\uu2.un19_w_addr_userZ0Z_0 ));
    CascadeMux I__2541 (
            .O(N__12345),
            .I(\uu2.un21_w_addr_displaying_i_cascade_ ));
    CascadeMux I__2540 (
            .O(N__12342),
            .I(N__12339));
    InMux I__2539 (
            .O(N__12339),
            .I(N__12334));
    InMux I__2538 (
            .O(N__12338),
            .I(N__12329));
    InMux I__2537 (
            .O(N__12337),
            .I(N__12329));
    LocalMux I__2536 (
            .O(N__12334),
            .I(\uu2.un15_w_data_displaying ));
    LocalMux I__2535 (
            .O(N__12329),
            .I(\uu2.un15_w_data_displaying ));
    InMux I__2534 (
            .O(N__12324),
            .I(N__12317));
    InMux I__2533 (
            .O(N__12323),
            .I(N__12317));
    CascadeMux I__2532 (
            .O(N__12322),
            .I(N__12312));
    LocalMux I__2531 (
            .O(N__12317),
            .I(N__12309));
    InMux I__2530 (
            .O(N__12316),
            .I(N__12306));
    CascadeMux I__2529 (
            .O(N__12315),
            .I(N__12302));
    InMux I__2528 (
            .O(N__12312),
            .I(N__12299));
    Span4Mux_h I__2527 (
            .O(N__12309),
            .I(N__12294));
    LocalMux I__2526 (
            .O(N__12306),
            .I(N__12294));
    CascadeMux I__2525 (
            .O(N__12305),
            .I(N__12288));
    InMux I__2524 (
            .O(N__12302),
            .I(N__12285));
    LocalMux I__2523 (
            .O(N__12299),
            .I(N__12282));
    Span4Mux_v I__2522 (
            .O(N__12294),
            .I(N__12279));
    InMux I__2521 (
            .O(N__12293),
            .I(N__12276));
    InMux I__2520 (
            .O(N__12292),
            .I(N__12269));
    InMux I__2519 (
            .O(N__12291),
            .I(N__12269));
    InMux I__2518 (
            .O(N__12288),
            .I(N__12269));
    LocalMux I__2517 (
            .O(N__12285),
            .I(N__12266));
    Span4Mux_h I__2516 (
            .O(N__12282),
            .I(N__12263));
    Odrv4 I__2515 (
            .O(N__12279),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2514 (
            .O(N__12276),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2513 (
            .O(N__12269),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv12 I__2512 (
            .O(N__12266),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__2511 (
            .O(N__12263),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    InMux I__2510 (
            .O(N__12252),
            .I(N__12249));
    LocalMux I__2509 (
            .O(N__12249),
            .I(\uu2.w_addr_displaying_4_0_i_rep1_6 ));
    CascadeMux I__2508 (
            .O(N__12246),
            .I(\uu2.w_addr_displaying_5_rep1_RNI3HMTZ0_cascade_ ));
    CascadeMux I__2507 (
            .O(N__12243),
            .I(\Lab_UT.didpuu0.countEnStens_cascade_ ));
    InMux I__2506 (
            .O(N__12240),
            .I(N__12237));
    LocalMux I__2505 (
            .O(N__12237),
            .I(\uu2.un1_segment4_2_amZ0Z_1 ));
    CascadeMux I__2504 (
            .O(N__12234),
            .I(\uu2.w_addr_displaying_4_0_i_6_cascade_ ));
    InMux I__2503 (
            .O(N__12231),
            .I(N__12226));
    InMux I__2502 (
            .O(N__12230),
            .I(N__12217));
    InMux I__2501 (
            .O(N__12229),
            .I(N__12217));
    LocalMux I__2500 (
            .O(N__12226),
            .I(N__12214));
    CascadeMux I__2499 (
            .O(N__12225),
            .I(N__12209));
    InMux I__2498 (
            .O(N__12224),
            .I(N__12204));
    InMux I__2497 (
            .O(N__12223),
            .I(N__12204));
    InMux I__2496 (
            .O(N__12222),
            .I(N__12201));
    LocalMux I__2495 (
            .O(N__12217),
            .I(N__12198));
    Span4Mux_v I__2494 (
            .O(N__12214),
            .I(N__12195));
    InMux I__2493 (
            .O(N__12213),
            .I(N__12192));
    InMux I__2492 (
            .O(N__12212),
            .I(N__12187));
    InMux I__2491 (
            .O(N__12209),
            .I(N__12187));
    LocalMux I__2490 (
            .O(N__12204),
            .I(N__12182));
    LocalMux I__2489 (
            .O(N__12201),
            .I(N__12182));
    Span4Mux_h I__2488 (
            .O(N__12198),
            .I(N__12178));
    Span4Mux_h I__2487 (
            .O(N__12195),
            .I(N__12173));
    LocalMux I__2486 (
            .O(N__12192),
            .I(N__12173));
    LocalMux I__2485 (
            .O(N__12187),
            .I(N__12168));
    Span4Mux_v I__2484 (
            .O(N__12182),
            .I(N__12168));
    InMux I__2483 (
            .O(N__12181),
            .I(N__12165));
    Odrv4 I__2482 (
            .O(N__12178),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2481 (
            .O(N__12173),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2480 (
            .O(N__12168),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2479 (
            .O(N__12165),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    CascadeMux I__2478 (
            .O(N__12156),
            .I(N__12153));
    InMux I__2477 (
            .O(N__12153),
            .I(N__12150));
    LocalMux I__2476 (
            .O(N__12150),
            .I(N__12147));
    Odrv4 I__2475 (
            .O(N__12147),
            .I(\uu2.g0_i_o4_0_a8_3_1 ));
    CascadeMux I__2474 (
            .O(N__12144),
            .I(uu2_un3_r_clk_en_0_cascade_));
    CascadeMux I__2473 (
            .O(N__12141),
            .I(N__12138));
    InMux I__2472 (
            .O(N__12138),
            .I(N__12135));
    LocalMux I__2471 (
            .O(N__12135),
            .I(\uu2.un349_ci_0 ));
    CascadeMux I__2470 (
            .O(N__12132),
            .I(N__12127));
    InMux I__2469 (
            .O(N__12131),
            .I(N__12124));
    InMux I__2468 (
            .O(N__12130),
            .I(N__12119));
    InMux I__2467 (
            .O(N__12127),
            .I(N__12119));
    LocalMux I__2466 (
            .O(N__12124),
            .I(\uu2.l_countZ0Z_7 ));
    LocalMux I__2465 (
            .O(N__12119),
            .I(\uu2.l_countZ0Z_7 ));
    InMux I__2464 (
            .O(N__12114),
            .I(N__12105));
    InMux I__2463 (
            .O(N__12113),
            .I(N__12105));
    InMux I__2462 (
            .O(N__12112),
            .I(N__12105));
    LocalMux I__2461 (
            .O(N__12105),
            .I(\uu2.l_countZ0Z_9 ));
    CascadeMux I__2460 (
            .O(N__12102),
            .I(N__12098));
    InMux I__2459 (
            .O(N__12101),
            .I(N__12094));
    InMux I__2458 (
            .O(N__12098),
            .I(N__12089));
    InMux I__2457 (
            .O(N__12097),
            .I(N__12089));
    LocalMux I__2456 (
            .O(N__12094),
            .I(N__12086));
    LocalMux I__2455 (
            .O(N__12089),
            .I(N__12083));
    Odrv4 I__2454 (
            .O(N__12086),
            .I(\uu2.vbuf_count.un382_ci_8_1 ));
    Odrv4 I__2453 (
            .O(N__12083),
            .I(\uu2.vbuf_count.un382_ci_8_1 ));
    CascadeMux I__2452 (
            .O(N__12078),
            .I(N__12072));
    InMux I__2451 (
            .O(N__12077),
            .I(N__12069));
    InMux I__2450 (
            .O(N__12076),
            .I(N__12064));
    InMux I__2449 (
            .O(N__12075),
            .I(N__12064));
    InMux I__2448 (
            .O(N__12072),
            .I(N__12061));
    LocalMux I__2447 (
            .O(N__12069),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__2446 (
            .O(N__12064),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__2445 (
            .O(N__12061),
            .I(\uu2.l_countZ0Z_8 ));
    CascadeMux I__2444 (
            .O(N__12054),
            .I(N__12049));
    InMux I__2443 (
            .O(N__12053),
            .I(N__12041));
    InMux I__2442 (
            .O(N__12052),
            .I(N__12041));
    InMux I__2441 (
            .O(N__12049),
            .I(N__12041));
    InMux I__2440 (
            .O(N__12048),
            .I(N__12036));
    LocalMux I__2439 (
            .O(N__12041),
            .I(N__12033));
    InMux I__2438 (
            .O(N__12040),
            .I(N__12028));
    InMux I__2437 (
            .O(N__12039),
            .I(N__12028));
    LocalMux I__2436 (
            .O(N__12036),
            .I(\uu2.l_countZ0Z_4 ));
    Odrv4 I__2435 (
            .O(N__12033),
            .I(\uu2.l_countZ0Z_4 ));
    LocalMux I__2434 (
            .O(N__12028),
            .I(\uu2.l_countZ0Z_4 ));
    CascadeMux I__2433 (
            .O(N__12021),
            .I(N__12018));
    InMux I__2432 (
            .O(N__12018),
            .I(N__12013));
    InMux I__2431 (
            .O(N__12017),
            .I(N__12010));
    CascadeMux I__2430 (
            .O(N__12016),
            .I(N__12003));
    LocalMux I__2429 (
            .O(N__12013),
            .I(N__11998));
    LocalMux I__2428 (
            .O(N__12010),
            .I(N__11998));
    InMux I__2427 (
            .O(N__12009),
            .I(N__11995));
    InMux I__2426 (
            .O(N__12008),
            .I(N__11986));
    InMux I__2425 (
            .O(N__12007),
            .I(N__11986));
    InMux I__2424 (
            .O(N__12006),
            .I(N__11986));
    InMux I__2423 (
            .O(N__12003),
            .I(N__11986));
    Odrv4 I__2422 (
            .O(N__11998),
            .I(\uu2.un316_ci ));
    LocalMux I__2421 (
            .O(N__11995),
            .I(\uu2.un316_ci ));
    LocalMux I__2420 (
            .O(N__11986),
            .I(\uu2.un316_ci ));
    InMux I__2419 (
            .O(N__11979),
            .I(N__11972));
    InMux I__2418 (
            .O(N__11978),
            .I(N__11967));
    InMux I__2417 (
            .O(N__11977),
            .I(N__11967));
    InMux I__2416 (
            .O(N__11976),
            .I(N__11962));
    InMux I__2415 (
            .O(N__11975),
            .I(N__11962));
    LocalMux I__2414 (
            .O(N__11972),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__2413 (
            .O(N__11967),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__2412 (
            .O(N__11962),
            .I(\uu2.l_countZ0Z_5 ));
    InMux I__2411 (
            .O(N__11955),
            .I(N__11949));
    InMux I__2410 (
            .O(N__11954),
            .I(N__11946));
    InMux I__2409 (
            .O(N__11953),
            .I(N__11943));
    InMux I__2408 (
            .O(N__11952),
            .I(N__11940));
    LocalMux I__2407 (
            .O(N__11949),
            .I(N__11937));
    LocalMux I__2406 (
            .O(N__11946),
            .I(\uu2.l_countZ0Z_6 ));
    LocalMux I__2405 (
            .O(N__11943),
            .I(\uu2.l_countZ0Z_6 ));
    LocalMux I__2404 (
            .O(N__11940),
            .I(\uu2.l_countZ0Z_6 ));
    Odrv4 I__2403 (
            .O(N__11937),
            .I(\uu2.l_countZ0Z_6 ));
    InMux I__2402 (
            .O(N__11928),
            .I(N__11925));
    LocalMux I__2401 (
            .O(N__11925),
            .I(\uu2.un382_ci ));
    InMux I__2400 (
            .O(N__11922),
            .I(N__11915));
    InMux I__2399 (
            .O(N__11921),
            .I(N__11910));
    InMux I__2398 (
            .O(N__11920),
            .I(N__11907));
    InMux I__2397 (
            .O(N__11919),
            .I(N__11904));
    InMux I__2396 (
            .O(N__11918),
            .I(N__11901));
    LocalMux I__2395 (
            .O(N__11915),
            .I(N__11898));
    InMux I__2394 (
            .O(N__11914),
            .I(N__11893));
    InMux I__2393 (
            .O(N__11913),
            .I(N__11893));
    LocalMux I__2392 (
            .O(N__11910),
            .I(uu2_un3_r_clk_en_0));
    LocalMux I__2391 (
            .O(N__11907),
            .I(uu2_un3_r_clk_en_0));
    LocalMux I__2390 (
            .O(N__11904),
            .I(uu2_un3_r_clk_en_0));
    LocalMux I__2389 (
            .O(N__11901),
            .I(uu2_un3_r_clk_en_0));
    Odrv4 I__2388 (
            .O(N__11898),
            .I(uu2_un3_r_clk_en_0));
    LocalMux I__2387 (
            .O(N__11893),
            .I(uu2_un3_r_clk_en_0));
    InMux I__2386 (
            .O(N__11880),
            .I(N__11876));
    InMux I__2385 (
            .O(N__11879),
            .I(N__11873));
    LocalMux I__2384 (
            .O(N__11876),
            .I(\uu2.l_countZ0Z_10 ));
    LocalMux I__2383 (
            .O(N__11873),
            .I(\uu2.l_countZ0Z_10 ));
    CascadeMux I__2382 (
            .O(N__11868),
            .I(\Lab_UT.didpuu0.countEnMones_cascade_ ));
    CEMux I__2381 (
            .O(N__11865),
            .I(N__11862));
    LocalMux I__2380 (
            .O(N__11862),
            .I(N__11859));
    Span4Mux_h I__2379 (
            .O(N__11859),
            .I(N__11856));
    Span4Mux_v I__2378 (
            .O(N__11856),
            .I(N__11853));
    Odrv4 I__2377 (
            .O(N__11853),
            .I(\Lab_UT.didpuu0.didpmones.countEnMones_0 ));
    CascadeMux I__2376 (
            .O(N__11850),
            .I(N__11845));
    CascadeMux I__2375 (
            .O(N__11849),
            .I(N__11842));
    InMux I__2374 (
            .O(N__11848),
            .I(N__11836));
    InMux I__2373 (
            .O(N__11845),
            .I(N__11836));
    InMux I__2372 (
            .O(N__11842),
            .I(N__11831));
    InMux I__2371 (
            .O(N__11841),
            .I(N__11831));
    LocalMux I__2370 (
            .O(N__11836),
            .I(\uu2.l_countZ0Z_2 ));
    LocalMux I__2369 (
            .O(N__11831),
            .I(\uu2.l_countZ0Z_2 ));
    InMux I__2368 (
            .O(N__11826),
            .I(N__11812));
    InMux I__2367 (
            .O(N__11825),
            .I(N__11812));
    InMux I__2366 (
            .O(N__11824),
            .I(N__11812));
    InMux I__2365 (
            .O(N__11823),
            .I(N__11812));
    InMux I__2364 (
            .O(N__11822),
            .I(N__11807));
    InMux I__2363 (
            .O(N__11821),
            .I(N__11807));
    LocalMux I__2362 (
            .O(N__11812),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__2361 (
            .O(N__11807),
            .I(\uu2.l_countZ0Z_0 ));
    CascadeMux I__2360 (
            .O(N__11802),
            .I(N__11799));
    InMux I__2359 (
            .O(N__11799),
            .I(N__11792));
    InMux I__2358 (
            .O(N__11798),
            .I(N__11792));
    InMux I__2357 (
            .O(N__11797),
            .I(N__11789));
    LocalMux I__2356 (
            .O(N__11792),
            .I(\uu2.l_countZ0Z_3 ));
    LocalMux I__2355 (
            .O(N__11789),
            .I(\uu2.l_countZ0Z_3 ));
    InMux I__2354 (
            .O(N__11784),
            .I(N__11771));
    InMux I__2353 (
            .O(N__11783),
            .I(N__11771));
    InMux I__2352 (
            .O(N__11782),
            .I(N__11771));
    InMux I__2351 (
            .O(N__11781),
            .I(N__11771));
    InMux I__2350 (
            .O(N__11780),
            .I(N__11768));
    LocalMux I__2349 (
            .O(N__11771),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__2348 (
            .O(N__11768),
            .I(\uu2.l_countZ0Z_1 ));
    InMux I__2347 (
            .O(N__11763),
            .I(N__11760));
    LocalMux I__2346 (
            .O(N__11760),
            .I(\uu2.un3_r_clk_en_7 ));
    CascadeMux I__2345 (
            .O(N__11757),
            .I(\uu2.un3_r_clk_en_0_0_cascade_ ));
    InMux I__2344 (
            .O(N__11754),
            .I(N__11751));
    LocalMux I__2343 (
            .O(N__11751),
            .I(\uu2.un3_r_clk_en_6 ));
    InMux I__2342 (
            .O(N__11748),
            .I(N__11745));
    LocalMux I__2341 (
            .O(N__11745),
            .I(N__11742));
    Span12Mux_s6_h I__2340 (
            .O(N__11742),
            .I(N__11739));
    Odrv12 I__2339 (
            .O(N__11739),
            .I(\uu2.mem0.G_14_0_a6_2_1 ));
    InMux I__2338 (
            .O(N__11736),
            .I(N__11733));
    LocalMux I__2337 (
            .O(N__11733),
            .I(\uu2.mem0.bitmap_pmux_1_1_2_tz_0 ));
    CascadeMux I__2336 (
            .O(N__11730),
            .I(N__11727));
    InMux I__2335 (
            .O(N__11727),
            .I(N__11724));
    LocalMux I__2334 (
            .O(N__11724),
            .I(\uu2.bitmap_pmux_1_1_2_tz_1_0 ));
    CascadeMux I__2333 (
            .O(N__11721),
            .I(\uu2.bitmap_pmux_1_1_2_tz_1_0_cascade_ ));
    CascadeMux I__2332 (
            .O(N__11718),
            .I(\uu2.mem0.bitmap_pmux_1_1_2_tz_cascade_ ));
    InMux I__2331 (
            .O(N__11715),
            .I(N__11712));
    LocalMux I__2330 (
            .O(N__11712),
            .I(N__11709));
    Span4Mux_v I__2329 (
            .O(N__11709),
            .I(N__11706));
    Odrv4 I__2328 (
            .O(N__11706),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_33 ));
    InMux I__2327 (
            .O(N__11703),
            .I(N__11700));
    LocalMux I__2326 (
            .O(N__11700),
            .I(N__11695));
    InMux I__2325 (
            .O(N__11699),
            .I(N__11691));
    InMux I__2324 (
            .O(N__11698),
            .I(N__11688));
    Span4Mux_h I__2323 (
            .O(N__11695),
            .I(N__11680));
    InMux I__2322 (
            .O(N__11694),
            .I(N__11677));
    LocalMux I__2321 (
            .O(N__11691),
            .I(N__11674));
    LocalMux I__2320 (
            .O(N__11688),
            .I(N__11671));
    InMux I__2319 (
            .O(N__11687),
            .I(N__11664));
    InMux I__2318 (
            .O(N__11686),
            .I(N__11664));
    InMux I__2317 (
            .O(N__11685),
            .I(N__11664));
    CascadeMux I__2316 (
            .O(N__11684),
            .I(N__11658));
    CascadeMux I__2315 (
            .O(N__11683),
            .I(N__11655));
    Span4Mux_v I__2314 (
            .O(N__11680),
            .I(N__11652));
    LocalMux I__2313 (
            .O(N__11677),
            .I(N__11649));
    Span4Mux_v I__2312 (
            .O(N__11674),
            .I(N__11642));
    Span4Mux_h I__2311 (
            .O(N__11671),
            .I(N__11642));
    LocalMux I__2310 (
            .O(N__11664),
            .I(N__11642));
    InMux I__2309 (
            .O(N__11663),
            .I(N__11631));
    InMux I__2308 (
            .O(N__11662),
            .I(N__11631));
    InMux I__2307 (
            .O(N__11661),
            .I(N__11631));
    InMux I__2306 (
            .O(N__11658),
            .I(N__11631));
    InMux I__2305 (
            .O(N__11655),
            .I(N__11631));
    Odrv4 I__2304 (
            .O(N__11652),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2303 (
            .O(N__11649),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2302 (
            .O(N__11642),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__2301 (
            .O(N__11631),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    CascadeMux I__2300 (
            .O(N__11622),
            .I(\uu2.w_addr_displaying_RNI8NHB1Z0Z_2_cascade_ ));
    InMux I__2299 (
            .O(N__11619),
            .I(N__11616));
    LocalMux I__2298 (
            .O(N__11616),
            .I(N__11613));
    Span4Mux_v I__2297 (
            .O(N__11613),
            .I(N__11610));
    Odrv4 I__2296 (
            .O(N__11610),
            .I(\uu2.w_addr_displaying_RNI18582Z0Z_8 ));
    CascadeMux I__2295 (
            .O(N__11607),
            .I(N__11603));
    CascadeMux I__2294 (
            .O(N__11606),
            .I(N__11600));
    InMux I__2293 (
            .O(N__11603),
            .I(N__11590));
    InMux I__2292 (
            .O(N__11600),
            .I(N__11590));
    CascadeMux I__2291 (
            .O(N__11599),
            .I(N__11583));
    InMux I__2290 (
            .O(N__11598),
            .I(N__11580));
    InMux I__2289 (
            .O(N__11597),
            .I(N__11575));
    InMux I__2288 (
            .O(N__11596),
            .I(N__11575));
    InMux I__2287 (
            .O(N__11595),
            .I(N__11572));
    LocalMux I__2286 (
            .O(N__11590),
            .I(N__11569));
    InMux I__2285 (
            .O(N__11589),
            .I(N__11562));
    InMux I__2284 (
            .O(N__11588),
            .I(N__11562));
    InMux I__2283 (
            .O(N__11587),
            .I(N__11562));
    InMux I__2282 (
            .O(N__11586),
            .I(N__11557));
    InMux I__2281 (
            .O(N__11583),
            .I(N__11557));
    LocalMux I__2280 (
            .O(N__11580),
            .I(\uu2.un1_w_addr_displaying_inv_4_0 ));
    LocalMux I__2279 (
            .O(N__11575),
            .I(\uu2.un1_w_addr_displaying_inv_4_0 ));
    LocalMux I__2278 (
            .O(N__11572),
            .I(\uu2.un1_w_addr_displaying_inv_4_0 ));
    Odrv4 I__2277 (
            .O(N__11569),
            .I(\uu2.un1_w_addr_displaying_inv_4_0 ));
    LocalMux I__2276 (
            .O(N__11562),
            .I(\uu2.un1_w_addr_displaying_inv_4_0 ));
    LocalMux I__2275 (
            .O(N__11557),
            .I(\uu2.un1_w_addr_displaying_inv_4_0 ));
    InMux I__2274 (
            .O(N__11544),
            .I(N__11541));
    LocalMux I__2273 (
            .O(N__11541),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_43 ));
    CascadeMux I__2272 (
            .O(N__11538),
            .I(\uu2.segment3_m_1Z0Z_6_cascade_ ));
    CascadeMux I__2271 (
            .O(N__11535),
            .I(\uu2.segment3_m_2_6_cascade_ ));
    InMux I__2270 (
            .O(N__11532),
            .I(N__11529));
    LocalMux I__2269 (
            .O(N__11529),
            .I(\uu2.un1_segment4_4_bmZ0 ));
    CascadeMux I__2268 (
            .O(N__11526),
            .I(\uu2.un1_segment4_4_amZ0_cascade_ ));
    CascadeMux I__2267 (
            .O(N__11523),
            .I(\uu2.N_111_cascade_ ));
    CascadeMux I__2266 (
            .O(N__11520),
            .I(\uu2.un1_segment4_sn_N_36_mux_0_cascade_ ));
    InMux I__2265 (
            .O(N__11517),
            .I(N__11514));
    LocalMux I__2264 (
            .O(N__11514),
            .I(N__11511));
    Odrv4 I__2263 (
            .O(N__11511),
            .I(\uu2.gZ0Z1 ));
    InMux I__2262 (
            .O(N__11508),
            .I(N__11505));
    LocalMux I__2261 (
            .O(N__11505),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_54 ));
    InMux I__2260 (
            .O(N__11502),
            .I(N__11499));
    LocalMux I__2259 (
            .O(N__11499),
            .I(\uu2.un1_segment4_sn_N_58_0 ));
    InMux I__2258 (
            .O(N__11496),
            .I(N__11493));
    LocalMux I__2257 (
            .O(N__11493),
            .I(\uu2.N_2150_0 ));
    InMux I__2256 (
            .O(N__11490),
            .I(N__11487));
    LocalMux I__2255 (
            .O(N__11487),
            .I(N__11484));
    Odrv4 I__2254 (
            .O(N__11484),
            .I(\uu2.un1_segment4_sn_N_38_0_0 ));
    CascadeMux I__2253 (
            .O(N__11481),
            .I(\uu2.g2_1_cascade_ ));
    InMux I__2252 (
            .O(N__11478),
            .I(N__11475));
    LocalMux I__2251 (
            .O(N__11475),
            .I(N__11472));
    Odrv4 I__2250 (
            .O(N__11472),
            .I(\uu2.N_299_0 ));
    CascadeMux I__2249 (
            .O(N__11469),
            .I(\uu2.g0_i_o4_0_a8_2_2_cascade_ ));
    InMux I__2248 (
            .O(N__11466),
            .I(N__11463));
    LocalMux I__2247 (
            .O(N__11463),
            .I(\uu2.w_addr_displaying_5_rep1_RNIVO2EZ0Z1 ));
    InMux I__2246 (
            .O(N__11460),
            .I(N__11457));
    LocalMux I__2245 (
            .O(N__11457),
            .I(N__11454));
    Odrv4 I__2244 (
            .O(N__11454),
            .I(\uu2.N_315_1_0 ));
    CascadeMux I__2243 (
            .O(N__11451),
            .I(N__11448));
    InMux I__2242 (
            .O(N__11448),
            .I(N__11445));
    LocalMux I__2241 (
            .O(N__11445),
            .I(\uu2.N_94 ));
    CascadeMux I__2240 (
            .O(N__11442),
            .I(\uu2.bitmap_pmux_1_1_3_tz_1_cascade_ ));
    InMux I__2239 (
            .O(N__11439),
            .I(N__11436));
    LocalMux I__2238 (
            .O(N__11436),
            .I(N__11432));
    InMux I__2237 (
            .O(N__11435),
            .I(N__11429));
    Span4Mux_h I__2236 (
            .O(N__11432),
            .I(N__11426));
    LocalMux I__2235 (
            .O(N__11429),
            .I(N__11423));
    Odrv4 I__2234 (
            .O(N__11426),
            .I(\uu2.bitmap_pmux_1_1_3_tz ));
    Odrv12 I__2233 (
            .O(N__11423),
            .I(\uu2.bitmap_pmux_1_1_3_tz ));
    CascadeMux I__2232 (
            .O(N__11418),
            .I(N__11415));
    InMux I__2231 (
            .O(N__11415),
            .I(N__11412));
    LocalMux I__2230 (
            .O(N__11412),
            .I(\Lab_UT.didpuu0.didpmtens.N_122 ));
    CascadeMux I__2229 (
            .O(N__11409),
            .I(N_84_cascade_));
    InMux I__2228 (
            .O(N__11406),
            .I(N__11402));
    InMux I__2227 (
            .O(N__11405),
            .I(N__11399));
    LocalMux I__2226 (
            .O(N__11402),
            .I(N_7));
    LocalMux I__2225 (
            .O(N__11399),
            .I(N_7));
    InMux I__2224 (
            .O(N__11394),
            .I(N__11391));
    LocalMux I__2223 (
            .O(N__11391),
            .I(\uu2.un1_segment4_0_bmZ0 ));
    CascadeMux I__2222 (
            .O(N__11388),
            .I(\uu2.un1_segment4_0_amZ0_cascade_ ));
    InMux I__2221 (
            .O(N__11385),
            .I(N__11382));
    LocalMux I__2220 (
            .O(N__11382),
            .I(N__11379));
    Span4Mux_v I__2219 (
            .O(N__11379),
            .I(N__11376));
    Odrv4 I__2218 (
            .O(N__11376),
            .I(\uu2.un1_segment4_2_bmZ0 ));
    CascadeMux I__2217 (
            .O(N__11373),
            .I(\uu2.un1_segment4_8_ns_1_cascade_ ));
    InMux I__2216 (
            .O(N__11370),
            .I(N__11367));
    LocalMux I__2215 (
            .O(N__11367),
            .I(\uu2.un1_segment4_2_amZ0 ));
    InMux I__2214 (
            .O(N__11364),
            .I(N__11361));
    LocalMux I__2213 (
            .O(N__11361),
            .I(\uu2.N_286 ));
    CascadeMux I__2212 (
            .O(N__11358),
            .I(\Lab_UT.N_10_cascade_ ));
    CascadeMux I__2211 (
            .O(N__11355),
            .I(vbuf_tx_data_rdy_cascade_));
    CEMux I__2210 (
            .O(N__11352),
            .I(N__11349));
    LocalMux I__2209 (
            .O(N__11349),
            .I(N__11345));
    CEMux I__2208 (
            .O(N__11348),
            .I(N__11342));
    Span4Mux_s3_h I__2207 (
            .O(N__11345),
            .I(N__11336));
    LocalMux I__2206 (
            .O(N__11342),
            .I(N__11336));
    CEMux I__2205 (
            .O(N__11341),
            .I(N__11333));
    Span4Mux_v I__2204 (
            .O(N__11336),
            .I(N__11328));
    LocalMux I__2203 (
            .O(N__11333),
            .I(N__11328));
    Span4Mux_h I__2202 (
            .O(N__11328),
            .I(N__11325));
    Odrv4 I__2201 (
            .O(N__11325),
            .I(\uu2.vbuf_tx_data_rdy_0 ));
    CascadeMux I__2200 (
            .O(N__11322),
            .I(N__11319));
    InMux I__2199 (
            .O(N__11319),
            .I(N__11316));
    LocalMux I__2198 (
            .O(N__11316),
            .I(N__11311));
    InMux I__2197 (
            .O(N__11315),
            .I(N__11306));
    InMux I__2196 (
            .O(N__11314),
            .I(N__11306));
    Span4Mux_v I__2195 (
            .O(N__11311),
            .I(N__11299));
    LocalMux I__2194 (
            .O(N__11306),
            .I(N__11299));
    InMux I__2193 (
            .O(N__11305),
            .I(N__11296));
    InMux I__2192 (
            .O(N__11304),
            .I(N__11293));
    Span4Mux_v I__2191 (
            .O(N__11299),
            .I(N__11290));
    LocalMux I__2190 (
            .O(N__11296),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__2189 (
            .O(N__11293),
            .I(\uu2.r_addrZ0Z_1 ));
    Odrv4 I__2188 (
            .O(N__11290),
            .I(\uu2.r_addrZ0Z_1 ));
    CascadeMux I__2187 (
            .O(N__11283),
            .I(N__11280));
    InMux I__2186 (
            .O(N__11280),
            .I(N__11276));
    InMux I__2185 (
            .O(N__11279),
            .I(N__11273));
    LocalMux I__2184 (
            .O(N__11276),
            .I(N__11269));
    LocalMux I__2183 (
            .O(N__11273),
            .I(N__11266));
    InMux I__2182 (
            .O(N__11272),
            .I(N__11263));
    Span4Mux_v I__2181 (
            .O(N__11269),
            .I(N__11256));
    Span4Mux_v I__2180 (
            .O(N__11266),
            .I(N__11256));
    LocalMux I__2179 (
            .O(N__11263),
            .I(N__11256));
    Span4Mux_h I__2178 (
            .O(N__11256),
            .I(N__11250));
    InMux I__2177 (
            .O(N__11255),
            .I(N__11247));
    InMux I__2176 (
            .O(N__11254),
            .I(N__11242));
    InMux I__2175 (
            .O(N__11253),
            .I(N__11242));
    Odrv4 I__2174 (
            .O(N__11250),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__2173 (
            .O(N__11247),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__2172 (
            .O(N__11242),
            .I(\uu2.r_addrZ0Z_0 ));
    CEMux I__2171 (
            .O(N__11235),
            .I(N__11229));
    InMux I__2170 (
            .O(N__11234),
            .I(N__11216));
    InMux I__2169 (
            .O(N__11233),
            .I(N__11216));
    SRMux I__2168 (
            .O(N__11232),
            .I(N__11213));
    LocalMux I__2167 (
            .O(N__11229),
            .I(N__11210));
    InMux I__2166 (
            .O(N__11228),
            .I(N__11193));
    InMux I__2165 (
            .O(N__11227),
            .I(N__11193));
    InMux I__2164 (
            .O(N__11226),
            .I(N__11193));
    InMux I__2163 (
            .O(N__11225),
            .I(N__11193));
    InMux I__2162 (
            .O(N__11224),
            .I(N__11193));
    InMux I__2161 (
            .O(N__11223),
            .I(N__11193));
    InMux I__2160 (
            .O(N__11222),
            .I(N__11193));
    InMux I__2159 (
            .O(N__11221),
            .I(N__11193));
    LocalMux I__2158 (
            .O(N__11216),
            .I(N__11186));
    LocalMux I__2157 (
            .O(N__11213),
            .I(N__11183));
    Span4Mux_v I__2156 (
            .O(N__11210),
            .I(N__11180));
    LocalMux I__2155 (
            .O(N__11193),
            .I(N__11177));
    InMux I__2154 (
            .O(N__11192),
            .I(N__11170));
    InMux I__2153 (
            .O(N__11191),
            .I(N__11170));
    InMux I__2152 (
            .O(N__11190),
            .I(N__11170));
    CascadeMux I__2151 (
            .O(N__11189),
            .I(N__11167));
    Span4Mux_h I__2150 (
            .O(N__11186),
            .I(N__11159));
    Span4Mux_v I__2149 (
            .O(N__11183),
            .I(N__11150));
    Span4Mux_s3_h I__2148 (
            .O(N__11180),
            .I(N__11150));
    Span4Mux_v I__2147 (
            .O(N__11177),
            .I(N__11150));
    LocalMux I__2146 (
            .O(N__11170),
            .I(N__11150));
    InMux I__2145 (
            .O(N__11167),
            .I(N__11147));
    InMux I__2144 (
            .O(N__11166),
            .I(N__11142));
    InMux I__2143 (
            .O(N__11165),
            .I(N__11142));
    InMux I__2142 (
            .O(N__11164),
            .I(N__11139));
    InMux I__2141 (
            .O(N__11163),
            .I(N__11136));
    InMux I__2140 (
            .O(N__11162),
            .I(N__11133));
    Span4Mux_v I__2139 (
            .O(N__11159),
            .I(N__11130));
    Span4Mux_v I__2138 (
            .O(N__11150),
            .I(N__11127));
    LocalMux I__2137 (
            .O(N__11147),
            .I(N__11120));
    LocalMux I__2136 (
            .O(N__11142),
            .I(N__11120));
    LocalMux I__2135 (
            .O(N__11139),
            .I(N__11120));
    LocalMux I__2134 (
            .O(N__11136),
            .I(vbuf_tx_data_rdy));
    LocalMux I__2133 (
            .O(N__11133),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__2132 (
            .O(N__11130),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__2131 (
            .O(N__11127),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__2130 (
            .O(N__11120),
            .I(vbuf_tx_data_rdy));
    CascadeMux I__2129 (
            .O(N__11109),
            .I(N__11106));
    InMux I__2128 (
            .O(N__11106),
            .I(N__11100));
    InMux I__2127 (
            .O(N__11105),
            .I(N__11095));
    InMux I__2126 (
            .O(N__11104),
            .I(N__11095));
    CascadeMux I__2125 (
            .O(N__11103),
            .I(N__11092));
    LocalMux I__2124 (
            .O(N__11100),
            .I(N__11087));
    LocalMux I__2123 (
            .O(N__11095),
            .I(N__11087));
    InMux I__2122 (
            .O(N__11092),
            .I(N__11084));
    Span4Mux_v I__2121 (
            .O(N__11087),
            .I(N__11081));
    LocalMux I__2120 (
            .O(N__11084),
            .I(\uu2.r_addrZ0Z_2 ));
    Odrv4 I__2119 (
            .O(N__11081),
            .I(\uu2.r_addrZ0Z_2 ));
    InMux I__2118 (
            .O(N__11076),
            .I(N__11073));
    LocalMux I__2117 (
            .O(N__11073),
            .I(N__11065));
    InMux I__2116 (
            .O(N__11072),
            .I(N__11058));
    InMux I__2115 (
            .O(N__11071),
            .I(N__11058));
    InMux I__2114 (
            .O(N__11070),
            .I(N__11058));
    InMux I__2113 (
            .O(N__11069),
            .I(N__11053));
    InMux I__2112 (
            .O(N__11068),
            .I(N__11053));
    Span4Mux_h I__2111 (
            .O(N__11065),
            .I(N__11049));
    LocalMux I__2110 (
            .O(N__11058),
            .I(N__11046));
    LocalMux I__2109 (
            .O(N__11053),
            .I(N__11037));
    InMux I__2108 (
            .O(N__11052),
            .I(N__11034));
    Span4Mux_h I__2107 (
            .O(N__11049),
            .I(N__11031));
    Span4Mux_h I__2106 (
            .O(N__11046),
            .I(N__11028));
    InMux I__2105 (
            .O(N__11045),
            .I(N__11025));
    InMux I__2104 (
            .O(N__11044),
            .I(N__11018));
    InMux I__2103 (
            .O(N__11043),
            .I(N__11018));
    InMux I__2102 (
            .O(N__11042),
            .I(N__11018));
    InMux I__2101 (
            .O(N__11041),
            .I(N__11013));
    InMux I__2100 (
            .O(N__11040),
            .I(N__11013));
    Span4Mux_h I__2099 (
            .O(N__11037),
            .I(N__11008));
    LocalMux I__2098 (
            .O(N__11034),
            .I(N__11008));
    Odrv4 I__2097 (
            .O(N__11031),
            .I(\Lab_UT.secuu0.un4_l_count_0 ));
    Odrv4 I__2096 (
            .O(N__11028),
            .I(\Lab_UT.secuu0.un4_l_count_0 ));
    LocalMux I__2095 (
            .O(N__11025),
            .I(\Lab_UT.secuu0.un4_l_count_0 ));
    LocalMux I__2094 (
            .O(N__11018),
            .I(\Lab_UT.secuu0.un4_l_count_0 ));
    LocalMux I__2093 (
            .O(N__11013),
            .I(\Lab_UT.secuu0.un4_l_count_0 ));
    Odrv4 I__2092 (
            .O(N__11008),
            .I(\Lab_UT.secuu0.un4_l_count_0 ));
    InMux I__2091 (
            .O(N__10995),
            .I(N__10992));
    LocalMux I__2090 (
            .O(N__10992),
            .I(N__10989));
    Span4Mux_h I__2089 (
            .O(N__10989),
            .I(N__10985));
    InMux I__2088 (
            .O(N__10988),
            .I(N__10982));
    Span4Mux_h I__2087 (
            .O(N__10985),
            .I(N__10977));
    LocalMux I__2086 (
            .O(N__10982),
            .I(N__10977));
    Odrv4 I__2085 (
            .O(N__10977),
            .I(\Lab_UT.secuu0.delay_lineZ0Z_0 ));
    InMux I__2084 (
            .O(N__10974),
            .I(N__10971));
    LocalMux I__2083 (
            .O(N__10971),
            .I(N__10968));
    Span4Mux_s3_h I__2082 (
            .O(N__10968),
            .I(N__10965));
    Odrv4 I__2081 (
            .O(N__10965),
            .I(\Lab_UT.secuu0.delay_lineZ0Z_1 ));
    InMux I__2080 (
            .O(N__10962),
            .I(N__10959));
    LocalMux I__2079 (
            .O(N__10959),
            .I(\resetGen.N_117 ));
    CascadeMux I__2078 (
            .O(N__10956),
            .I(N__10952));
    InMux I__2077 (
            .O(N__10955),
            .I(N__10949));
    InMux I__2076 (
            .O(N__10952),
            .I(N__10946));
    LocalMux I__2075 (
            .O(N__10949),
            .I(\resetGen.reset_countZ0Z_3 ));
    LocalMux I__2074 (
            .O(N__10946),
            .I(\resetGen.reset_countZ0Z_3 ));
    CascadeMux I__2073 (
            .O(N__10941),
            .I(\resetGen.N_117_cascade_ ));
    InMux I__2072 (
            .O(N__10938),
            .I(N__10935));
    LocalMux I__2071 (
            .O(N__10935),
            .I(N__10932));
    Span4Mux_v I__2070 (
            .O(N__10932),
            .I(N__10928));
    IoInMux I__2069 (
            .O(N__10931),
            .I(N__10925));
    IoSpan4Mux I__2068 (
            .O(N__10928),
            .I(N__10920));
    LocalMux I__2067 (
            .O(N__10925),
            .I(N__10920));
    IoSpan4Mux I__2066 (
            .O(N__10920),
            .I(N__10917));
    Span4Mux_s3_h I__2065 (
            .O(N__10917),
            .I(N__10914));
    Odrv4 I__2064 (
            .O(N__10914),
            .I(rst));
    CascadeMux I__2063 (
            .O(N__10911),
            .I(N__10908));
    InMux I__2062 (
            .O(N__10908),
            .I(N__10896));
    InMux I__2061 (
            .O(N__10907),
            .I(N__10896));
    InMux I__2060 (
            .O(N__10906),
            .I(N__10896));
    InMux I__2059 (
            .O(N__10905),
            .I(N__10896));
    LocalMux I__2058 (
            .O(N__10896),
            .I(\resetGen.reset_countZ0Z_0 ));
    InMux I__2057 (
            .O(N__10893),
            .I(N__10884));
    InMux I__2056 (
            .O(N__10892),
            .I(N__10884));
    InMux I__2055 (
            .O(N__10891),
            .I(N__10884));
    LocalMux I__2054 (
            .O(N__10884),
            .I(\resetGen.reset_countZ0Z_1 ));
    InMux I__2053 (
            .O(N__10881),
            .I(N__10873));
    InMux I__2052 (
            .O(N__10880),
            .I(N__10868));
    InMux I__2051 (
            .O(N__10879),
            .I(N__10868));
    InMux I__2050 (
            .O(N__10878),
            .I(N__10861));
    InMux I__2049 (
            .O(N__10877),
            .I(N__10861));
    InMux I__2048 (
            .O(N__10876),
            .I(N__10861));
    LocalMux I__2047 (
            .O(N__10873),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__2046 (
            .O(N__10868),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__2045 (
            .O(N__10861),
            .I(\resetGen.reset_countZ0Z_4 ));
    CascadeMux I__2044 (
            .O(N__10854),
            .I(\resetGen.N_96_cascade_ ));
    InMux I__2043 (
            .O(N__10851),
            .I(N__10839));
    InMux I__2042 (
            .O(N__10850),
            .I(N__10839));
    InMux I__2041 (
            .O(N__10849),
            .I(N__10839));
    InMux I__2040 (
            .O(N__10848),
            .I(N__10839));
    LocalMux I__2039 (
            .O(N__10839),
            .I(N__10835));
    InMux I__2038 (
            .O(N__10838),
            .I(N__10832));
    Span4Mux_h I__2037 (
            .O(N__10835),
            .I(N__10829));
    LocalMux I__2036 (
            .O(N__10832),
            .I(\resetGen.N_133 ));
    Odrv4 I__2035 (
            .O(N__10829),
            .I(\resetGen.N_133 ));
    InMux I__2034 (
            .O(N__10824),
            .I(N__10818));
    InMux I__2033 (
            .O(N__10823),
            .I(N__10818));
    LocalMux I__2032 (
            .O(N__10818),
            .I(\resetGen.reset_countZ0Z_2 ));
    InMux I__2031 (
            .O(N__10815),
            .I(N__10808));
    InMux I__2030 (
            .O(N__10814),
            .I(N__10805));
    CascadeMux I__2029 (
            .O(N__10813),
            .I(N__10802));
    InMux I__2028 (
            .O(N__10812),
            .I(N__10798));
    InMux I__2027 (
            .O(N__10811),
            .I(N__10795));
    LocalMux I__2026 (
            .O(N__10808),
            .I(N__10790));
    LocalMux I__2025 (
            .O(N__10805),
            .I(N__10790));
    InMux I__2024 (
            .O(N__10802),
            .I(N__10785));
    InMux I__2023 (
            .O(N__10801),
            .I(N__10785));
    LocalMux I__2022 (
            .O(N__10798),
            .I(buart__tx_uart_busy_0));
    LocalMux I__2021 (
            .O(N__10795),
            .I(buart__tx_uart_busy_0));
    Odrv4 I__2020 (
            .O(N__10790),
            .I(buart__tx_uart_busy_0));
    LocalMux I__2019 (
            .O(N__10785),
            .I(buart__tx_uart_busy_0));
    InMux I__2018 (
            .O(N__10776),
            .I(\buart.Z_tx.un1_bitcount_cry_0 ));
    InMux I__2017 (
            .O(N__10773),
            .I(\buart.Z_tx.un1_bitcount_cry_1 ));
    InMux I__2016 (
            .O(N__10770),
            .I(N__10767));
    LocalMux I__2015 (
            .O(N__10767),
            .I(\buart.Z_tx.un1_bitcount_axb_3 ));
    InMux I__2014 (
            .O(N__10764),
            .I(\buart.Z_tx.un1_bitcount_cry_2 ));
    InMux I__2013 (
            .O(N__10761),
            .I(N__10758));
    LocalMux I__2012 (
            .O(N__10758),
            .I(\buart.Z_tx.bitcount_RNIM5O32Z0Z_2 ));
    InMux I__2011 (
            .O(N__10755),
            .I(N__10752));
    LocalMux I__2010 (
            .O(N__10752),
            .I(\buart.Z_tx.bitcount_RNIL4O32Z0Z_1 ));
    CascadeMux I__2009 (
            .O(N__10749),
            .I(N__10745));
    InMux I__2008 (
            .O(N__10748),
            .I(N__10741));
    InMux I__2007 (
            .O(N__10745),
            .I(N__10736));
    InMux I__2006 (
            .O(N__10744),
            .I(N__10736));
    LocalMux I__2005 (
            .O(N__10741),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    LocalMux I__2004 (
            .O(N__10736),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__2003 (
            .O(N__10731),
            .I(N__10727));
    InMux I__2002 (
            .O(N__10730),
            .I(N__10719));
    InMux I__2001 (
            .O(N__10727),
            .I(N__10719));
    InMux I__2000 (
            .O(N__10726),
            .I(N__10719));
    LocalMux I__1999 (
            .O(N__10719),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    CascadeMux I__1998 (
            .O(N__10716),
            .I(N__10712));
    InMux I__1997 (
            .O(N__10715),
            .I(N__10709));
    InMux I__1996 (
            .O(N__10712),
            .I(N__10706));
    LocalMux I__1995 (
            .O(N__10709),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    LocalMux I__1994 (
            .O(N__10706),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    CascadeMux I__1993 (
            .O(N__10701),
            .I(N__10697));
    InMux I__1992 (
            .O(N__10700),
            .I(N__10692));
    InMux I__1991 (
            .O(N__10697),
            .I(N__10689));
    InMux I__1990 (
            .O(N__10696),
            .I(N__10684));
    InMux I__1989 (
            .O(N__10695),
            .I(N__10684));
    LocalMux I__1988 (
            .O(N__10692),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__1987 (
            .O(N__10689),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__1986 (
            .O(N__10684),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    CascadeMux I__1985 (
            .O(N__10677),
            .I(buart__tx_uart_busy_0_cascade_));
    InMux I__1984 (
            .O(N__10674),
            .I(N__10663));
    InMux I__1983 (
            .O(N__10673),
            .I(N__10656));
    InMux I__1982 (
            .O(N__10672),
            .I(N__10656));
    InMux I__1981 (
            .O(N__10671),
            .I(N__10656));
    InMux I__1980 (
            .O(N__10670),
            .I(N__10651));
    InMux I__1979 (
            .O(N__10669),
            .I(N__10651));
    InMux I__1978 (
            .O(N__10668),
            .I(N__10644));
    InMux I__1977 (
            .O(N__10667),
            .I(N__10644));
    InMux I__1976 (
            .O(N__10666),
            .I(N__10644));
    LocalMux I__1975 (
            .O(N__10663),
            .I(N__10641));
    LocalMux I__1974 (
            .O(N__10656),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__1973 (
            .O(N__10651),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__1972 (
            .O(N__10644),
            .I(\buart.Z_tx.ser_clk ));
    Odrv4 I__1971 (
            .O(N__10641),
            .I(\buart.Z_tx.ser_clk ));
    InMux I__1970 (
            .O(N__10632),
            .I(N__10629));
    LocalMux I__1969 (
            .O(N__10629),
            .I(\buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0 ));
    CascadeMux I__1968 (
            .O(N__10626),
            .I(N__10623));
    InMux I__1967 (
            .O(N__10623),
            .I(N__10620));
    LocalMux I__1966 (
            .O(N__10620),
            .I(N__10617));
    Odrv4 I__1965 (
            .O(N__10617),
            .I(\uu2.un1_segment4_5_bmZ0 ));
    CascadeMux I__1964 (
            .O(N__10614),
            .I(\Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMUZ0Z_0_cascade_ ));
    IoInMux I__1963 (
            .O(N__10611),
            .I(N__10608));
    LocalMux I__1962 (
            .O(N__10608),
            .I(N__10605));
    Span4Mux_s2_h I__1961 (
            .O(N__10605),
            .I(N__10602));
    Span4Mux_h I__1960 (
            .O(N__10602),
            .I(N__10599));
    Odrv4 I__1959 (
            .O(N__10599),
            .I(led_c_2));
    InMux I__1958 (
            .O(N__10596),
            .I(N__10593));
    LocalMux I__1957 (
            .O(N__10593),
            .I(\Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJZ0Z_0 ));
    InMux I__1956 (
            .O(N__10590),
            .I(N__10587));
    LocalMux I__1955 (
            .O(N__10587),
            .I(N__10584));
    Odrv4 I__1954 (
            .O(N__10584),
            .I(\uu2.un1_segment4_5_amZ0Z_1 ));
    InMux I__1953 (
            .O(N__10581),
            .I(N__10578));
    LocalMux I__1952 (
            .O(N__10578),
            .I(\uu2.w_addr_displaying_fast_RNIV5694Z0Z_2 ));
    CascadeMux I__1951 (
            .O(N__10575),
            .I(\uu2.N_290_0_i_0_cascade_ ));
    InMux I__1950 (
            .O(N__10572),
            .I(N__10569));
    LocalMux I__1949 (
            .O(N__10569),
            .I(\uu2.w_addr_displaying_RNI362A1Z0Z_3 ));
    CascadeMux I__1948 (
            .O(N__10566),
            .I(\uu2.un1_w_addr_displaying_19_cascade_ ));
    CascadeMux I__1947 (
            .O(N__10563),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_ ));
    InMux I__1946 (
            .O(N__10560),
            .I(N__10557));
    LocalMux I__1945 (
            .O(N__10557),
            .I(N__10554));
    Span4Mux_h I__1944 (
            .O(N__10554),
            .I(N__10551));
    Odrv4 I__1943 (
            .O(N__10551),
            .I(\uu2.mem0.N_5_0 ));
    InMux I__1942 (
            .O(N__10548),
            .I(N__10543));
    InMux I__1941 (
            .O(N__10547),
            .I(N__10540));
    InMux I__1940 (
            .O(N__10546),
            .I(N__10537));
    LocalMux I__1939 (
            .O(N__10543),
            .I(N__10532));
    LocalMux I__1938 (
            .O(N__10540),
            .I(N__10532));
    LocalMux I__1937 (
            .O(N__10537),
            .I(\uu2.un1_segment3_s_0 ));
    Odrv4 I__1936 (
            .O(N__10532),
            .I(\uu2.un1_segment3_s_0 ));
    InMux I__1935 (
            .O(N__10527),
            .I(N__10523));
    InMux I__1934 (
            .O(N__10526),
            .I(N__10520));
    LocalMux I__1933 (
            .O(N__10523),
            .I(\uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4 ));
    LocalMux I__1932 (
            .O(N__10520),
            .I(\uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4 ));
    InMux I__1931 (
            .O(N__10515),
            .I(N__10512));
    LocalMux I__1930 (
            .O(N__10512),
            .I(\uu2.mem0.un1_segment3_m2_2 ));
    InMux I__1929 (
            .O(N__10509),
            .I(N__10506));
    LocalMux I__1928 (
            .O(N__10506),
            .I(\uu2.mem0.un1_segment3_m2_0 ));
    CascadeMux I__1927 (
            .O(N__10503),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_42_cascade_ ));
    InMux I__1926 (
            .O(N__10500),
            .I(N__10497));
    LocalMux I__1925 (
            .O(N__10497),
            .I(N__10494));
    Odrv4 I__1924 (
            .O(N__10494),
            .I(\uu2.mem0.un1_segment3_1_0 ));
    InMux I__1923 (
            .O(N__10491),
            .I(N__10488));
    LocalMux I__1922 (
            .O(N__10488),
            .I(N__10485));
    Span4Mux_v I__1921 (
            .O(N__10485),
            .I(N__10482));
    Odrv4 I__1920 (
            .O(N__10482),
            .I(\Lab_UT.didpuu0.didpmtens.q_5_0_0_2 ));
    InMux I__1919 (
            .O(N__10479),
            .I(N__10476));
    LocalMux I__1918 (
            .O(N__10476),
            .I(N__10473));
    Odrv12 I__1917 (
            .O(N__10473),
            .I(\uu2.un1_segment4_1_amZ0 ));
    CascadeMux I__1916 (
            .O(N__10470),
            .I(\uu2.un1_segment4_1_bmZ0_cascade_ ));
    CascadeMux I__1915 (
            .O(N__10467),
            .I(\uu2.w_addr_displaying_fast_RNIPN54Z0Z_8_cascade_ ));
    InMux I__1914 (
            .O(N__10464),
            .I(N__10461));
    LocalMux I__1913 (
            .O(N__10461),
            .I(N__10458));
    Odrv4 I__1912 (
            .O(N__10458),
            .I(\uu2.N_292 ));
    InMux I__1911 (
            .O(N__10455),
            .I(N__10451));
    InMux I__1910 (
            .O(N__10454),
            .I(N__10448));
    LocalMux I__1909 (
            .O(N__10451),
            .I(\uu2.N_93 ));
    LocalMux I__1908 (
            .O(N__10448),
            .I(\uu2.N_93 ));
    CascadeMux I__1907 (
            .O(N__10443),
            .I(\uu2.N_49_cascade_ ));
    InMux I__1906 (
            .O(N__10440),
            .I(N__10437));
    LocalMux I__1905 (
            .O(N__10437),
            .I(\uu2.un1_segment3_m4_s_2 ));
    InMux I__1904 (
            .O(N__10434),
            .I(N__10431));
    LocalMux I__1903 (
            .O(N__10431),
            .I(\uu2.g0_i_o4_0_1 ));
    InMux I__1902 (
            .O(N__10428),
            .I(N__10425));
    LocalMux I__1901 (
            .O(N__10425),
            .I(\uu2.un1_segment3_m4_ns_1 ));
    CascadeMux I__1900 (
            .O(N__10422),
            .I(\uu2.g0_i_o4_3_cascade_ ));
    InMux I__1899 (
            .O(N__10419),
            .I(N__10415));
    CascadeMux I__1898 (
            .O(N__10418),
            .I(N__10410));
    LocalMux I__1897 (
            .O(N__10415),
            .I(N__10407));
    InMux I__1896 (
            .O(N__10414),
            .I(N__10400));
    InMux I__1895 (
            .O(N__10413),
            .I(N__10400));
    InMux I__1894 (
            .O(N__10410),
            .I(N__10400));
    Odrv4 I__1893 (
            .O(N__10407),
            .I(\uu2.un1_segment3_m4 ));
    LocalMux I__1892 (
            .O(N__10400),
            .I(\uu2.un1_segment3_m4 ));
    InMux I__1891 (
            .O(N__10395),
            .I(N__10392));
    LocalMux I__1890 (
            .O(N__10392),
            .I(\uu2.w_addr_displaying_4_rep1_RNIMMRIAZ0 ));
    CascadeMux I__1889 (
            .O(N__10389),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_53_cascade_ ));
    InMux I__1888 (
            .O(N__10386),
            .I(N__10383));
    LocalMux I__1887 (
            .O(N__10383),
            .I(\uu2.mem0.un1_segment3_1_2 ));
    CascadeMux I__1886 (
            .O(N__10380),
            .I(Lab_UT_dec3_segmentUQ_1_1_cascade_));
    InMux I__1885 (
            .O(N__10377),
            .I(N__10374));
    LocalMux I__1884 (
            .O(N__10374),
            .I(\uu2.Z_decfrac105_7_2 ));
    InMux I__1883 (
            .O(N__10371),
            .I(N__10366));
    CascadeMux I__1882 (
            .O(N__10370),
            .I(N__10361));
    CascadeMux I__1881 (
            .O(N__10369),
            .I(N__10358));
    LocalMux I__1880 (
            .O(N__10366),
            .I(N__10355));
    InMux I__1879 (
            .O(N__10365),
            .I(N__10350));
    InMux I__1878 (
            .O(N__10364),
            .I(N__10350));
    InMux I__1877 (
            .O(N__10361),
            .I(N__10347));
    InMux I__1876 (
            .O(N__10358),
            .I(N__10344));
    Span4Mux_v I__1875 (
            .O(N__10355),
            .I(N__10339));
    LocalMux I__1874 (
            .O(N__10350),
            .I(N__10339));
    LocalMux I__1873 (
            .O(N__10347),
            .I(N__10336));
    LocalMux I__1872 (
            .O(N__10344),
            .I(N__10333));
    Span4Mux_h I__1871 (
            .O(N__10339),
            .I(N__10330));
    Span4Mux_v I__1870 (
            .O(N__10336),
            .I(N__10325));
    Span4Mux_v I__1869 (
            .O(N__10333),
            .I(N__10325));
    Odrv4 I__1868 (
            .O(N__10330),
            .I(\Lab_UT.rx_data_0 ));
    Odrv4 I__1867 (
            .O(N__10325),
            .I(\Lab_UT.rx_data_0 ));
    CascadeMux I__1866 (
            .O(N__10320),
            .I(N__10317));
    InMux I__1865 (
            .O(N__10317),
            .I(N__10313));
    InMux I__1864 (
            .O(N__10316),
            .I(N__10309));
    LocalMux I__1863 (
            .O(N__10313),
            .I(N__10306));
    InMux I__1862 (
            .O(N__10312),
            .I(N__10303));
    LocalMux I__1861 (
            .O(N__10309),
            .I(N__10298));
    Span4Mux_v I__1860 (
            .O(N__10306),
            .I(N__10298));
    LocalMux I__1859 (
            .O(N__10303),
            .I(N__10294));
    Span4Mux_h I__1858 (
            .O(N__10298),
            .I(N__10291));
    InMux I__1857 (
            .O(N__10297),
            .I(N__10288));
    Odrv12 I__1856 (
            .O(N__10294),
            .I(\Lab_UT.rx_dataZ0Z_2 ));
    Odrv4 I__1855 (
            .O(N__10291),
            .I(\Lab_UT.rx_dataZ0Z_2 ));
    LocalMux I__1854 (
            .O(N__10288),
            .I(\Lab_UT.rx_dataZ0Z_2 ));
    InMux I__1853 (
            .O(N__10281),
            .I(N__10278));
    LocalMux I__1852 (
            .O(N__10278),
            .I(\Lab_UT.dictrluu0.N_103_1 ));
    InMux I__1851 (
            .O(N__10275),
            .I(N__10272));
    LocalMux I__1850 (
            .O(N__10272),
            .I(N__10269));
    Odrv4 I__1849 (
            .O(N__10269),
            .I(\Lab_UT.dicSelectLEDdisp ));
    CascadeMux I__1848 (
            .O(N__10266),
            .I(\Lab_UT.dicSelectLEDdisp_cascade_ ));
    InMux I__1847 (
            .O(N__10263),
            .I(N__10257));
    InMux I__1846 (
            .O(N__10262),
            .I(N__10257));
    LocalMux I__1845 (
            .O(N__10257),
            .I(N__10254));
    Odrv4 I__1844 (
            .O(N__10254),
            .I(\Lab_UT.dictrluu0.N_72 ));
    InMux I__1843 (
            .O(N__10251),
            .I(N__10248));
    LocalMux I__1842 (
            .O(N__10248),
            .I(\Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_o2_2 ));
    InMux I__1841 (
            .O(N__10245),
            .I(N__10242));
    LocalMux I__1840 (
            .O(N__10242),
            .I(N__10239));
    Odrv4 I__1839 (
            .O(N__10239),
            .I(\Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_3 ));
    InMux I__1838 (
            .O(N__10236),
            .I(N__10233));
    LocalMux I__1837 (
            .O(N__10233),
            .I(\Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_4 ));
    CascadeMux I__1836 (
            .O(N__10230),
            .I(\Lab_UT.dictrluu0.dicfsm.N_102_cascade_ ));
    InMux I__1835 (
            .O(N__10227),
            .I(N__10219));
    InMux I__1834 (
            .O(N__10226),
            .I(N__10219));
    CascadeMux I__1833 (
            .O(N__10225),
            .I(N__10216));
    CascadeMux I__1832 (
            .O(N__10224),
            .I(N__10213));
    LocalMux I__1831 (
            .O(N__10219),
            .I(N__10210));
    InMux I__1830 (
            .O(N__10216),
            .I(N__10207));
    InMux I__1829 (
            .O(N__10213),
            .I(N__10204));
    Odrv12 I__1828 (
            .O(N__10210),
            .I(Lab_UT_rx_data_7));
    LocalMux I__1827 (
            .O(N__10207),
            .I(Lab_UT_rx_data_7));
    LocalMux I__1826 (
            .O(N__10204),
            .I(Lab_UT_rx_data_7));
    InMux I__1825 (
            .O(N__10197),
            .I(N__10192));
    InMux I__1824 (
            .O(N__10196),
            .I(N__10187));
    InMux I__1823 (
            .O(N__10195),
            .I(N__10187));
    LocalMux I__1822 (
            .O(N__10192),
            .I(N__10184));
    LocalMux I__1821 (
            .O(N__10187),
            .I(N__10179));
    Span4Mux_s3_h I__1820 (
            .O(N__10184),
            .I(N__10176));
    InMux I__1819 (
            .O(N__10183),
            .I(N__10171));
    InMux I__1818 (
            .O(N__10182),
            .I(N__10171));
    Odrv4 I__1817 (
            .O(N__10179),
            .I(Lab_UT_rx_data_1));
    Odrv4 I__1816 (
            .O(N__10176),
            .I(Lab_UT_rx_data_1));
    LocalMux I__1815 (
            .O(N__10171),
            .I(Lab_UT_rx_data_1));
    CascadeMux I__1814 (
            .O(N__10164),
            .I(N__10160));
    CascadeMux I__1813 (
            .O(N__10163),
            .I(N__10156));
    InMux I__1812 (
            .O(N__10160),
            .I(N__10150));
    InMux I__1811 (
            .O(N__10159),
            .I(N__10150));
    InMux I__1810 (
            .O(N__10156),
            .I(N__10147));
    CascadeMux I__1809 (
            .O(N__10155),
            .I(N__10144));
    LocalMux I__1808 (
            .O(N__10150),
            .I(N__10141));
    LocalMux I__1807 (
            .O(N__10147),
            .I(N__10138));
    InMux I__1806 (
            .O(N__10144),
            .I(N__10135));
    Odrv12 I__1805 (
            .O(N__10141),
            .I(Lab_UT_rx_data_6));
    Odrv4 I__1804 (
            .O(N__10138),
            .I(Lab_UT_rx_data_6));
    LocalMux I__1803 (
            .O(N__10135),
            .I(Lab_UT_rx_data_6));
    CascadeMux I__1802 (
            .O(N__10128),
            .I(N__10124));
    InMux I__1801 (
            .O(N__10127),
            .I(N__10119));
    InMux I__1800 (
            .O(N__10124),
            .I(N__10119));
    LocalMux I__1799 (
            .O(N__10119),
            .I(\Lab_UT.rx_data_rdy ));
    InMux I__1798 (
            .O(N__10116),
            .I(N__10106));
    InMux I__1797 (
            .O(N__10115),
            .I(N__10106));
    InMux I__1796 (
            .O(N__10114),
            .I(N__10100));
    InMux I__1795 (
            .O(N__10113),
            .I(N__10100));
    InMux I__1794 (
            .O(N__10112),
            .I(N__10097));
    InMux I__1793 (
            .O(N__10111),
            .I(N__10094));
    LocalMux I__1792 (
            .O(N__10106),
            .I(N__10091));
    InMux I__1791 (
            .O(N__10105),
            .I(N__10088));
    LocalMux I__1790 (
            .O(N__10100),
            .I(N__10085));
    LocalMux I__1789 (
            .O(N__10097),
            .I(buart__rx_bitcount_0));
    LocalMux I__1788 (
            .O(N__10094),
            .I(buart__rx_bitcount_0));
    Odrv4 I__1787 (
            .O(N__10091),
            .I(buart__rx_bitcount_0));
    LocalMux I__1786 (
            .O(N__10088),
            .I(buart__rx_bitcount_0));
    Odrv4 I__1785 (
            .O(N__10085),
            .I(buart__rx_bitcount_0));
    InMux I__1784 (
            .O(N__10074),
            .I(N__10064));
    InMux I__1783 (
            .O(N__10073),
            .I(N__10064));
    InMux I__1782 (
            .O(N__10072),
            .I(N__10060));
    InMux I__1781 (
            .O(N__10071),
            .I(N__10055));
    InMux I__1780 (
            .O(N__10070),
            .I(N__10055));
    InMux I__1779 (
            .O(N__10069),
            .I(N__10052));
    LocalMux I__1778 (
            .O(N__10064),
            .I(N__10049));
    InMux I__1777 (
            .O(N__10063),
            .I(N__10046));
    LocalMux I__1776 (
            .O(N__10060),
            .I(N__10043));
    LocalMux I__1775 (
            .O(N__10055),
            .I(buart__rx_bitcount_2));
    LocalMux I__1774 (
            .O(N__10052),
            .I(buart__rx_bitcount_2));
    Odrv4 I__1773 (
            .O(N__10049),
            .I(buart__rx_bitcount_2));
    LocalMux I__1772 (
            .O(N__10046),
            .I(buart__rx_bitcount_2));
    Odrv4 I__1771 (
            .O(N__10043),
            .I(buart__rx_bitcount_2));
    CascadeMux I__1770 (
            .O(N__10032),
            .I(N__10027));
    CascadeMux I__1769 (
            .O(N__10031),
            .I(N__10024));
    CascadeMux I__1768 (
            .O(N__10030),
            .I(N__10020));
    InMux I__1767 (
            .O(N__10027),
            .I(N__10015));
    InMux I__1766 (
            .O(N__10024),
            .I(N__10015));
    CascadeMux I__1765 (
            .O(N__10023),
            .I(N__10010));
    InMux I__1764 (
            .O(N__10020),
            .I(N__10006));
    LocalMux I__1763 (
            .O(N__10015),
            .I(N__10003));
    InMux I__1762 (
            .O(N__10014),
            .I(N__10000));
    InMux I__1761 (
            .O(N__10013),
            .I(N__9997));
    InMux I__1760 (
            .O(N__10010),
            .I(N__9994));
    InMux I__1759 (
            .O(N__10009),
            .I(N__9991));
    LocalMux I__1758 (
            .O(N__10006),
            .I(N__9988));
    Span4Mux_h I__1757 (
            .O(N__10003),
            .I(N__9985));
    LocalMux I__1756 (
            .O(N__10000),
            .I(buart__rx_bitcount_3));
    LocalMux I__1755 (
            .O(N__9997),
            .I(buart__rx_bitcount_3));
    LocalMux I__1754 (
            .O(N__9994),
            .I(buart__rx_bitcount_3));
    LocalMux I__1753 (
            .O(N__9991),
            .I(buart__rx_bitcount_3));
    Odrv4 I__1752 (
            .O(N__9988),
            .I(buart__rx_bitcount_3));
    Odrv4 I__1751 (
            .O(N__9985),
            .I(buart__rx_bitcount_3));
    InMux I__1750 (
            .O(N__9972),
            .I(N__9964));
    InMux I__1749 (
            .O(N__9971),
            .I(N__9964));
    InMux I__1748 (
            .O(N__9970),
            .I(N__9961));
    InMux I__1747 (
            .O(N__9969),
            .I(N__9958));
    LocalMux I__1746 (
            .O(N__9964),
            .I(N__9955));
    LocalMux I__1745 (
            .O(N__9961),
            .I(N__9952));
    LocalMux I__1744 (
            .O(N__9958),
            .I(N_118));
    Odrv4 I__1743 (
            .O(N__9955),
            .I(N_118));
    Odrv4 I__1742 (
            .O(N__9952),
            .I(N_118));
    InMux I__1741 (
            .O(N__9945),
            .I(N__9939));
    InMux I__1740 (
            .O(N__9944),
            .I(N__9939));
    LocalMux I__1739 (
            .O(N__9939),
            .I(bu_rx_data_rdy));
    InMux I__1738 (
            .O(N__9936),
            .I(N__9931));
    InMux I__1737 (
            .O(N__9935),
            .I(N__9925));
    InMux I__1736 (
            .O(N__9934),
            .I(N__9925));
    LocalMux I__1735 (
            .O(N__9931),
            .I(N__9922));
    InMux I__1734 (
            .O(N__9930),
            .I(N__9919));
    LocalMux I__1733 (
            .O(N__9925),
            .I(\buart.Z_rx.ser_clk ));
    Odrv12 I__1732 (
            .O(N__9922),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__1731 (
            .O(N__9919),
            .I(\buart.Z_rx.ser_clk ));
    InMux I__1730 (
            .O(N__9912),
            .I(N__9908));
    InMux I__1729 (
            .O(N__9911),
            .I(N__9905));
    LocalMux I__1728 (
            .O(N__9908),
            .I(\buart.Z_rx.N_129 ));
    LocalMux I__1727 (
            .O(N__9905),
            .I(\buart.Z_rx.N_129 ));
    CascadeMux I__1726 (
            .O(N__9900),
            .I(bu_rx_data_rdy_cascade_));
    CascadeMux I__1725 (
            .O(N__9897),
            .I(N__9893));
    CascadeMux I__1724 (
            .O(N__9896),
            .I(N__9890));
    InMux I__1723 (
            .O(N__9893),
            .I(N__9885));
    InMux I__1722 (
            .O(N__9890),
            .I(N__9880));
    InMux I__1721 (
            .O(N__9889),
            .I(N__9880));
    CascadeMux I__1720 (
            .O(N__9888),
            .I(N__9876));
    LocalMux I__1719 (
            .O(N__9885),
            .I(N__9865));
    LocalMux I__1718 (
            .O(N__9880),
            .I(N__9865));
    InMux I__1717 (
            .O(N__9879),
            .I(N__9862));
    InMux I__1716 (
            .O(N__9876),
            .I(N__9853));
    InMux I__1715 (
            .O(N__9875),
            .I(N__9853));
    InMux I__1714 (
            .O(N__9874),
            .I(N__9853));
    InMux I__1713 (
            .O(N__9873),
            .I(N__9853));
    InMux I__1712 (
            .O(N__9872),
            .I(N__9846));
    InMux I__1711 (
            .O(N__9871),
            .I(N__9846));
    InMux I__1710 (
            .O(N__9870),
            .I(N__9846));
    Span4Mux_s3_v I__1709 (
            .O(N__9865),
            .I(N__9842));
    LocalMux I__1708 (
            .O(N__9862),
            .I(N__9835));
    LocalMux I__1707 (
            .O(N__9853),
            .I(N__9835));
    LocalMux I__1706 (
            .O(N__9846),
            .I(N__9835));
    InMux I__1705 (
            .O(N__9845),
            .I(N__9832));
    Odrv4 I__1704 (
            .O(N__9842),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__1703 (
            .O(N__9835),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__1702 (
            .O(N__9832),
            .I(\buart.Z_rx.startbit ));
    CEMux I__1701 (
            .O(N__9825),
            .I(N__9821));
    CEMux I__1700 (
            .O(N__9824),
            .I(N__9818));
    LocalMux I__1699 (
            .O(N__9821),
            .I(N__9815));
    LocalMux I__1698 (
            .O(N__9818),
            .I(N__9812));
    Span4Mux_s3_v I__1697 (
            .O(N__9815),
            .I(N__9807));
    Span4Mux_h I__1696 (
            .O(N__9812),
            .I(N__9807));
    Odrv4 I__1695 (
            .O(N__9807),
            .I(\buart.Z_rx.bitcount_e_0_RNII0231Z0Z_0 ));
    CascadeMux I__1694 (
            .O(N__9804),
            .I(Lab_UT_dec3_segmentUQ_0_6_cascade_));
    InMux I__1693 (
            .O(N__9801),
            .I(N__9798));
    LocalMux I__1692 (
            .O(N__9798),
            .I(N_71));
    CascadeMux I__1691 (
            .O(N__9795),
            .I(N_71_cascade_));
    InMux I__1690 (
            .O(N__9792),
            .I(N__9785));
    InMux I__1689 (
            .O(N__9791),
            .I(N__9785));
    InMux I__1688 (
            .O(N__9790),
            .I(N__9782));
    LocalMux I__1687 (
            .O(N__9785),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__1686 (
            .O(N__9782),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    InMux I__1685 (
            .O(N__9777),
            .I(N__9773));
    InMux I__1684 (
            .O(N__9776),
            .I(N__9770));
    LocalMux I__1683 (
            .O(N__9773),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    LocalMux I__1682 (
            .O(N__9770),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__1681 (
            .O(N__9765),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ));
    CascadeMux I__1680 (
            .O(N__9762),
            .I(N__9756));
    InMux I__1679 (
            .O(N__9761),
            .I(N__9749));
    InMux I__1678 (
            .O(N__9760),
            .I(N__9749));
    InMux I__1677 (
            .O(N__9759),
            .I(N__9749));
    InMux I__1676 (
            .O(N__9756),
            .I(N__9746));
    LocalMux I__1675 (
            .O(N__9749),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1674 (
            .O(N__9746),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__1673 (
            .O(N__9741),
            .I(N__9738));
    LocalMux I__1672 (
            .O(N__9738),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    CascadeMux I__1671 (
            .O(N__9735),
            .I(\buart.Z_rx.ser_clk_cascade_ ));
    InMux I__1670 (
            .O(N__9732),
            .I(N__9727));
    InMux I__1669 (
            .O(N__9731),
            .I(N__9722));
    InMux I__1668 (
            .O(N__9730),
            .I(N__9722));
    LocalMux I__1667 (
            .O(N__9727),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__1666 (
            .O(N__9722),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    InMux I__1665 (
            .O(N__9717),
            .I(N__9714));
    LocalMux I__1664 (
            .O(N__9714),
            .I(N__9710));
    InMux I__1663 (
            .O(N__9713),
            .I(N__9706));
    Span4Mux_h I__1662 (
            .O(N__9710),
            .I(N__9703));
    InMux I__1661 (
            .O(N__9709),
            .I(N__9700));
    LocalMux I__1660 (
            .O(N__9706),
            .I(N__9697));
    Odrv4 I__1659 (
            .O(N__9703),
            .I(bu_rx_data_7));
    LocalMux I__1658 (
            .O(N__9700),
            .I(bu_rx_data_7));
    Odrv4 I__1657 (
            .O(N__9697),
            .I(bu_rx_data_7));
    InMux I__1656 (
            .O(N__9690),
            .I(N__9687));
    LocalMux I__1655 (
            .O(N__9687),
            .I(N__9683));
    CascadeMux I__1654 (
            .O(N__9686),
            .I(N__9679));
    Span4Mux_h I__1653 (
            .O(N__9683),
            .I(N__9676));
    InMux I__1652 (
            .O(N__9682),
            .I(N__9671));
    InMux I__1651 (
            .O(N__9679),
            .I(N__9671));
    Odrv4 I__1650 (
            .O(N__9676),
            .I(bu_rx_data_6));
    LocalMux I__1649 (
            .O(N__9671),
            .I(bu_rx_data_6));
    InMux I__1648 (
            .O(N__9666),
            .I(N__9663));
    LocalMux I__1647 (
            .O(N__9663),
            .I(N__9660));
    Span12Mux_s5_h I__1646 (
            .O(N__9660),
            .I(N__9655));
    InMux I__1645 (
            .O(N__9659),
            .I(N__9652));
    InMux I__1644 (
            .O(N__9658),
            .I(N__9649));
    Odrv12 I__1643 (
            .O(N__9655),
            .I(bu_rx_data_2));
    LocalMux I__1642 (
            .O(N__9652),
            .I(bu_rx_data_2));
    LocalMux I__1641 (
            .O(N__9649),
            .I(bu_rx_data_2));
    InMux I__1640 (
            .O(N__9642),
            .I(N__9639));
    LocalMux I__1639 (
            .O(N__9639),
            .I(N__9636));
    Span4Mux_h I__1638 (
            .O(N__9636),
            .I(N__9631));
    InMux I__1637 (
            .O(N__9635),
            .I(N__9628));
    InMux I__1636 (
            .O(N__9634),
            .I(N__9625));
    Odrv4 I__1635 (
            .O(N__9631),
            .I(bu_rx_data_4));
    LocalMux I__1634 (
            .O(N__9628),
            .I(bu_rx_data_4));
    LocalMux I__1633 (
            .O(N__9625),
            .I(bu_rx_data_4));
    InMux I__1632 (
            .O(N__9618),
            .I(N__9615));
    LocalMux I__1631 (
            .O(N__9615),
            .I(N__9611));
    CascadeMux I__1630 (
            .O(N__9614),
            .I(N__9607));
    Span4Mux_v I__1629 (
            .O(N__9611),
            .I(N__9604));
    InMux I__1628 (
            .O(N__9610),
            .I(N__9601));
    InMux I__1627 (
            .O(N__9607),
            .I(N__9598));
    Odrv4 I__1626 (
            .O(N__9604),
            .I(bu_rx_data_3));
    LocalMux I__1625 (
            .O(N__9601),
            .I(bu_rx_data_3));
    LocalMux I__1624 (
            .O(N__9598),
            .I(bu_rx_data_3));
    InMux I__1623 (
            .O(N__9591),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__1622 (
            .O(N__9588),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__1621 (
            .O(N__9585),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    InMux I__1620 (
            .O(N__9582),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    CascadeMux I__1619 (
            .O(N__9579),
            .I(N__9576));
    InMux I__1618 (
            .O(N__9576),
            .I(N__9573));
    LocalMux I__1617 (
            .O(N__9573),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    CEMux I__1616 (
            .O(N__9570),
            .I(N__9567));
    LocalMux I__1615 (
            .O(N__9567),
            .I(N__9564));
    Span4Mux_v I__1614 (
            .O(N__9564),
            .I(N__9561));
    Span4Mux_s0_v I__1613 (
            .O(N__9561),
            .I(N__9557));
    CEMux I__1612 (
            .O(N__9560),
            .I(N__9554));
    Span4Mux_v I__1611 (
            .O(N__9557),
            .I(N__9549));
    LocalMux I__1610 (
            .O(N__9554),
            .I(N__9549));
    Span4Mux_v I__1609 (
            .O(N__9549),
            .I(N__9546));
    Span4Mux_v I__1608 (
            .O(N__9546),
            .I(N__9543));
    Odrv4 I__1607 (
            .O(N__9543),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    InMux I__1606 (
            .O(N__9540),
            .I(N__9536));
    InMux I__1605 (
            .O(N__9539),
            .I(N__9533));
    LocalMux I__1604 (
            .O(N__9536),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__1603 (
            .O(N__9533),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    CascadeMux I__1602 (
            .O(N__9528),
            .I(N__9523));
    InMux I__1601 (
            .O(N__9527),
            .I(N__9520));
    InMux I__1600 (
            .O(N__9526),
            .I(N__9515));
    InMux I__1599 (
            .O(N__9523),
            .I(N__9515));
    LocalMux I__1598 (
            .O(N__9520),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1597 (
            .O(N__9515),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    InMux I__1596 (
            .O(N__9510),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__1595 (
            .O(N__9507),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__1594 (
            .O(N__9504),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    CascadeMux I__1593 (
            .O(N__9501),
            .I(N__9498));
    InMux I__1592 (
            .O(N__9498),
            .I(N__9492));
    InMux I__1591 (
            .O(N__9497),
            .I(N__9492));
    LocalMux I__1590 (
            .O(N__9492),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__1589 (
            .O(N__9489),
            .I(N__9486));
    InMux I__1588 (
            .O(N__9486),
            .I(N__9480));
    InMux I__1587 (
            .O(N__9485),
            .I(N__9480));
    LocalMux I__1586 (
            .O(N__9480),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__1585 (
            .O(N__9477),
            .I(N__9473));
    InMux I__1584 (
            .O(N__9476),
            .I(N__9470));
    InMux I__1583 (
            .O(N__9473),
            .I(N__9467));
    LocalMux I__1582 (
            .O(N__9470),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    LocalMux I__1581 (
            .O(N__9467),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    CascadeMux I__1580 (
            .O(N__9462),
            .I(N__9459));
    InMux I__1579 (
            .O(N__9459),
            .I(N__9453));
    InMux I__1578 (
            .O(N__9458),
            .I(N__9453));
    LocalMux I__1577 (
            .O(N__9453),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    CascadeMux I__1576 (
            .O(N__9450),
            .I(N__9446));
    InMux I__1575 (
            .O(N__9449),
            .I(N__9441));
    InMux I__1574 (
            .O(N__9446),
            .I(N__9441));
    LocalMux I__1573 (
            .O(N__9441),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__1572 (
            .O(N__9438),
            .I(N__9435));
    LocalMux I__1571 (
            .O(N__9435),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    InMux I__1570 (
            .O(N__9432),
            .I(N__9424));
    InMux I__1569 (
            .O(N__9431),
            .I(N__9424));
    InMux I__1568 (
            .O(N__9430),
            .I(N__9421));
    InMux I__1567 (
            .O(N__9429),
            .I(N__9418));
    LocalMux I__1566 (
            .O(N__9424),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1565 (
            .O(N__9421),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1564 (
            .O(N__9418),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__1563 (
            .O(N__9411),
            .I(N__9407));
    InMux I__1562 (
            .O(N__9410),
            .I(N__9403));
    InMux I__1561 (
            .O(N__9407),
            .I(N__9400));
    InMux I__1560 (
            .O(N__9406),
            .I(N__9397));
    LocalMux I__1559 (
            .O(N__9403),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1558 (
            .O(N__9400),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1557 (
            .O(N__9397),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    InMux I__1556 (
            .O(N__9390),
            .I(N__9387));
    LocalMux I__1555 (
            .O(N__9387),
            .I(vbuf_tx_data_7));
    InMux I__1554 (
            .O(N__9384),
            .I(N__9381));
    LocalMux I__1553 (
            .O(N__9381),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CascadeMux I__1552 (
            .O(N__9378),
            .I(N__9375));
    InMux I__1551 (
            .O(N__9375),
            .I(N__9372));
    LocalMux I__1550 (
            .O(N__9372),
            .I(N__9367));
    InMux I__1549 (
            .O(N__9371),
            .I(N__9362));
    InMux I__1548 (
            .O(N__9370),
            .I(N__9359));
    Span4Mux_h I__1547 (
            .O(N__9367),
            .I(N__9356));
    InMux I__1546 (
            .O(N__9366),
            .I(N__9351));
    InMux I__1545 (
            .O(N__9365),
            .I(N__9351));
    LocalMux I__1544 (
            .O(N__9362),
            .I(\uu2.w_addr_userZ0Z_4 ));
    LocalMux I__1543 (
            .O(N__9359),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv4 I__1542 (
            .O(N__9356),
            .I(\uu2.w_addr_userZ0Z_4 ));
    LocalMux I__1541 (
            .O(N__9351),
            .I(\uu2.w_addr_userZ0Z_4 ));
    CascadeMux I__1540 (
            .O(N__9342),
            .I(N__9339));
    InMux I__1539 (
            .O(N__9339),
            .I(N__9336));
    LocalMux I__1538 (
            .O(N__9336),
            .I(N__9333));
    Span4Mux_h I__1537 (
            .O(N__9333),
            .I(N__9330));
    Odrv4 I__1536 (
            .O(N__9330),
            .I(\uu2.mem0.w_addr_4 ));
    InMux I__1535 (
            .O(N__9327),
            .I(N__9324));
    LocalMux I__1534 (
            .O(N__9324),
            .I(N__9319));
    CascadeMux I__1533 (
            .O(N__9323),
            .I(N__9315));
    InMux I__1532 (
            .O(N__9322),
            .I(N__9312));
    Span4Mux_h I__1531 (
            .O(N__9319),
            .I(N__9309));
    InMux I__1530 (
            .O(N__9318),
            .I(N__9304));
    InMux I__1529 (
            .O(N__9315),
            .I(N__9304));
    LocalMux I__1528 (
            .O(N__9312),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__1527 (
            .O(N__9309),
            .I(\uu2.w_addr_userZ0Z_5 ));
    LocalMux I__1526 (
            .O(N__9304),
            .I(\uu2.w_addr_userZ0Z_5 ));
    CascadeMux I__1525 (
            .O(N__9297),
            .I(N__9294));
    InMux I__1524 (
            .O(N__9294),
            .I(N__9291));
    LocalMux I__1523 (
            .O(N__9291),
            .I(N__9288));
    Span4Mux_v I__1522 (
            .O(N__9288),
            .I(N__9285));
    Span4Mux_s2_h I__1521 (
            .O(N__9285),
            .I(N__9282));
    Odrv4 I__1520 (
            .O(N__9282),
            .I(\uu2.mem0.w_addr_5 ));
    CascadeMux I__1519 (
            .O(N__9279),
            .I(N__9276));
    InMux I__1518 (
            .O(N__9276),
            .I(N__9273));
    LocalMux I__1517 (
            .O(N__9273),
            .I(N__9270));
    Odrv4 I__1516 (
            .O(N__9270),
            .I(\uu2.Z_decfrac106_2 ));
    InMux I__1515 (
            .O(N__9267),
            .I(N__9264));
    LocalMux I__1514 (
            .O(N__9264),
            .I(N__9261));
    Span4Mux_h I__1513 (
            .O(N__9261),
            .I(N__9258));
    Odrv4 I__1512 (
            .O(N__9258),
            .I(\uu2.mem0.N_2160_1 ));
    InMux I__1511 (
            .O(N__9255),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__1510 (
            .O(N__9252),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__1509 (
            .O(N__9249),
            .I(N__9246));
    LocalMux I__1508 (
            .O(N__9246),
            .I(\uu2.mem0.un1_segment3_0 ));
    InMux I__1507 (
            .O(N__9243),
            .I(N__9240));
    LocalMux I__1506 (
            .O(N__9240),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_34 ));
    CascadeMux I__1505 (
            .O(N__9237),
            .I(N__9232));
    CascadeMux I__1504 (
            .O(N__9236),
            .I(N__9229));
    InMux I__1503 (
            .O(N__9235),
            .I(N__9221));
    InMux I__1502 (
            .O(N__9232),
            .I(N__9221));
    InMux I__1501 (
            .O(N__9229),
            .I(N__9221));
    InMux I__1500 (
            .O(N__9228),
            .I(N__9218));
    LocalMux I__1499 (
            .O(N__9221),
            .I(N__9212));
    LocalMux I__1498 (
            .O(N__9218),
            .I(N__9212));
    InMux I__1497 (
            .O(N__9217),
            .I(N__9209));
    Odrv4 I__1496 (
            .O(N__9212),
            .I(\uu2.Z_decfrac106 ));
    LocalMux I__1495 (
            .O(N__9209),
            .I(\uu2.Z_decfrac106 ));
    InMux I__1494 (
            .O(N__9204),
            .I(N__9201));
    LocalMux I__1493 (
            .O(N__9201),
            .I(\uu2.mem0.un1_segment3_m2_1 ));
    CascadeMux I__1492 (
            .O(N__9198),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_47_cascade_ ));
    CascadeMux I__1491 (
            .O(N__9195),
            .I(N__9192));
    InMux I__1490 (
            .O(N__9192),
            .I(N__9189));
    LocalMux I__1489 (
            .O(N__9189),
            .I(\uu2.mem0.un1_segment3_1_1 ));
    InMux I__1488 (
            .O(N__9186),
            .I(N__9183));
    LocalMux I__1487 (
            .O(N__9183),
            .I(\uu2.mem0.N_2160_0 ));
    InMux I__1486 (
            .O(N__9180),
            .I(N__9177));
    LocalMux I__1485 (
            .O(N__9177),
            .I(N__9174));
    Odrv4 I__1484 (
            .O(N__9174),
            .I(N_52));
    InMux I__1483 (
            .O(N__9171),
            .I(N__9168));
    LocalMux I__1482 (
            .O(N__9168),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_48 ));
    InMux I__1481 (
            .O(N__9165),
            .I(N__9162));
    LocalMux I__1480 (
            .O(N__9162),
            .I(vbuf_tx_data_6));
    InMux I__1479 (
            .O(N__9159),
            .I(N__9156));
    LocalMux I__1478 (
            .O(N__9156),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__1477 (
            .O(N__9153),
            .I(N__9150));
    LocalMux I__1476 (
            .O(N__9150),
            .I(N__9147));
    Odrv4 I__1475 (
            .O(N__9147),
            .I(N_52_0));
    InMux I__1474 (
            .O(N__9144),
            .I(N__9141));
    LocalMux I__1473 (
            .O(N__9141),
            .I(L3_segment2_0_0));
    CascadeMux I__1472 (
            .O(N__9138),
            .I(\uu2.mem0.N_2159_0_cascade_ ));
    InMux I__1471 (
            .O(N__9135),
            .I(N__9132));
    LocalMux I__1470 (
            .O(N__9132),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_20 ));
    InMux I__1469 (
            .O(N__9129),
            .I(N__9126));
    LocalMux I__1468 (
            .O(N__9126),
            .I(N__9123));
    Odrv12 I__1467 (
            .O(N__9123),
            .I(L3_segment2_0));
    CascadeMux I__1466 (
            .O(N__9120),
            .I(\uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4_cascade_ ));
    InMux I__1465 (
            .O(N__9117),
            .I(N__9114));
    LocalMux I__1464 (
            .O(N__9114),
            .I(\uu2.mem0.g2_0 ));
    CascadeMux I__1463 (
            .O(N__9111),
            .I(\uu2.mem0.N_5_cascade_ ));
    InMux I__1462 (
            .O(N__9108),
            .I(N__9105));
    LocalMux I__1461 (
            .O(N__9105),
            .I(\uu2.mem0.bitmap_pmux_1_1_0_0 ));
    InMux I__1460 (
            .O(N__9102),
            .I(N__9099));
    LocalMux I__1459 (
            .O(N__9099),
            .I(\uu2.mem0.N_14 ));
    InMux I__1458 (
            .O(N__9096),
            .I(N__9093));
    LocalMux I__1457 (
            .O(N__9093),
            .I(\uu2.mem0.N_18 ));
    CEMux I__1456 (
            .O(N__9090),
            .I(N__9087));
    LocalMux I__1455 (
            .O(N__9087),
            .I(N__9084));
    Span4Mux_s1_h I__1454 (
            .O(N__9084),
            .I(N__9079));
    CEMux I__1453 (
            .O(N__9083),
            .I(N__9076));
    CEMux I__1452 (
            .O(N__9082),
            .I(N__9073));
    Span4Mux_v I__1451 (
            .O(N__9079),
            .I(N__9070));
    LocalMux I__1450 (
            .O(N__9076),
            .I(N__9067));
    LocalMux I__1449 (
            .O(N__9073),
            .I(N__9064));
    Span4Mux_h I__1448 (
            .O(N__9070),
            .I(N__9061));
    Span4Mux_s2_h I__1447 (
            .O(N__9067),
            .I(N__9058));
    Span4Mux_h I__1446 (
            .O(N__9064),
            .I(N__9055));
    Odrv4 I__1445 (
            .O(N__9061),
            .I(\Lab_UT.Lab3U00.bu_rx_data_rdy_0 ));
    Odrv4 I__1444 (
            .O(N__9058),
            .I(\Lab_UT.Lab3U00.bu_rx_data_rdy_0 ));
    Odrv4 I__1443 (
            .O(N__9055),
            .I(\Lab_UT.Lab3U00.bu_rx_data_rdy_0 ));
    InMux I__1442 (
            .O(N__9048),
            .I(N__9043));
    CascadeMux I__1441 (
            .O(N__9047),
            .I(N__9040));
    CascadeMux I__1440 (
            .O(N__9046),
            .I(N__9037));
    LocalMux I__1439 (
            .O(N__9043),
            .I(N__9032));
    InMux I__1438 (
            .O(N__9040),
            .I(N__9029));
    InMux I__1437 (
            .O(N__9037),
            .I(N__9026));
    InMux I__1436 (
            .O(N__9036),
            .I(N__9021));
    InMux I__1435 (
            .O(N__9035),
            .I(N__9021));
    Span4Mux_h I__1434 (
            .O(N__9032),
            .I(N__9018));
    LocalMux I__1433 (
            .O(N__9029),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__1432 (
            .O(N__9026),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__1431 (
            .O(N__9021),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv4 I__1430 (
            .O(N__9018),
            .I(\uu2.w_addr_userZ0Z_2 ));
    CascadeMux I__1429 (
            .O(N__9009),
            .I(N__9006));
    InMux I__1428 (
            .O(N__9006),
            .I(N__9003));
    LocalMux I__1427 (
            .O(N__9003),
            .I(N__9000));
    Span4Mux_v I__1426 (
            .O(N__9000),
            .I(N__8997));
    Odrv4 I__1425 (
            .O(N__8997),
            .I(\uu2.mem0.w_addr_2 ));
    InMux I__1424 (
            .O(N__8994),
            .I(N__8991));
    LocalMux I__1423 (
            .O(N__8991),
            .I(N__8984));
    InMux I__1422 (
            .O(N__8990),
            .I(N__8979));
    InMux I__1421 (
            .O(N__8989),
            .I(N__8979));
    InMux I__1420 (
            .O(N__8988),
            .I(N__8974));
    InMux I__1419 (
            .O(N__8987),
            .I(N__8974));
    Span4Mux_h I__1418 (
            .O(N__8984),
            .I(N__8971));
    LocalMux I__1417 (
            .O(N__8979),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__1416 (
            .O(N__8974),
            .I(\uu2.w_addr_userZ0Z_3 ));
    Odrv4 I__1415 (
            .O(N__8971),
            .I(\uu2.w_addr_userZ0Z_3 ));
    CascadeMux I__1414 (
            .O(N__8964),
            .I(N__8961));
    InMux I__1413 (
            .O(N__8961),
            .I(N__8958));
    LocalMux I__1412 (
            .O(N__8958),
            .I(N__8955));
    Span4Mux_h I__1411 (
            .O(N__8955),
            .I(N__8952));
    Odrv4 I__1410 (
            .O(N__8952),
            .I(\uu2.mem0.w_addr_3 ));
    InMux I__1409 (
            .O(N__8949),
            .I(N__8946));
    LocalMux I__1408 (
            .O(N__8946),
            .I(\uu2.mem0.G_14_0_0 ));
    CascadeMux I__1407 (
            .O(N__8943),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_32_cascade_ ));
    InMux I__1406 (
            .O(N__8940),
            .I(N__8937));
    LocalMux I__1405 (
            .O(N__8937),
            .I(\uu2.mem0.G_14_0_1 ));
    CascadeMux I__1404 (
            .O(N__8934),
            .I(\uu2.N_329_0_cascade_ ));
    CascadeMux I__1403 (
            .O(N__8931),
            .I(N__8928));
    InMux I__1402 (
            .O(N__8928),
            .I(N__8923));
    InMux I__1401 (
            .O(N__8927),
            .I(N__8920));
    InMux I__1400 (
            .O(N__8926),
            .I(N__8914));
    LocalMux I__1399 (
            .O(N__8923),
            .I(N__8911));
    LocalMux I__1398 (
            .O(N__8920),
            .I(N__8908));
    InMux I__1397 (
            .O(N__8919),
            .I(N__8903));
    InMux I__1396 (
            .O(N__8918),
            .I(N__8903));
    InMux I__1395 (
            .O(N__8917),
            .I(N__8900));
    LocalMux I__1394 (
            .O(N__8914),
            .I(N__8897));
    Odrv4 I__1393 (
            .O(N__8911),
            .I(\uu2.Z_decfrac105_7 ));
    Odrv4 I__1392 (
            .O(N__8908),
            .I(\uu2.Z_decfrac105_7 ));
    LocalMux I__1391 (
            .O(N__8903),
            .I(\uu2.Z_decfrac105_7 ));
    LocalMux I__1390 (
            .O(N__8900),
            .I(\uu2.Z_decfrac105_7 ));
    Odrv4 I__1389 (
            .O(N__8897),
            .I(\uu2.Z_decfrac105_7 ));
    CascadeMux I__1388 (
            .O(N__8886),
            .I(N__8882));
    InMux I__1387 (
            .O(N__8885),
            .I(N__8876));
    InMux I__1386 (
            .O(N__8882),
            .I(N__8867));
    InMux I__1385 (
            .O(N__8881),
            .I(N__8867));
    InMux I__1384 (
            .O(N__8880),
            .I(N__8867));
    InMux I__1383 (
            .O(N__8879),
            .I(N__8867));
    LocalMux I__1382 (
            .O(N__8876),
            .I(N__8862));
    LocalMux I__1381 (
            .O(N__8867),
            .I(N__8862));
    Odrv12 I__1380 (
            .O(N__8862),
            .I(\buart.Z_rx.N_39 ));
    CascadeMux I__1379 (
            .O(N__8859),
            .I(N__8854));
    InMux I__1378 (
            .O(N__8858),
            .I(N__8849));
    InMux I__1377 (
            .O(N__8857),
            .I(N__8849));
    InMux I__1376 (
            .O(N__8854),
            .I(N__8846));
    LocalMux I__1375 (
            .O(N__8849),
            .I(N__8843));
    LocalMux I__1374 (
            .O(N__8846),
            .I(N__8838));
    Span4Mux_v I__1373 (
            .O(N__8843),
            .I(N__8835));
    InMux I__1372 (
            .O(N__8842),
            .I(N__8832));
    InMux I__1371 (
            .O(N__8841),
            .I(N__8829));
    Odrv12 I__1370 (
            .O(N__8838),
            .I(Lab_UT_rx_data_4));
    Odrv4 I__1369 (
            .O(N__8835),
            .I(Lab_UT_rx_data_4));
    LocalMux I__1368 (
            .O(N__8832),
            .I(Lab_UT_rx_data_4));
    LocalMux I__1367 (
            .O(N__8829),
            .I(Lab_UT_rx_data_4));
    CascadeMux I__1366 (
            .O(N__8820),
            .I(N__8817));
    InMux I__1365 (
            .O(N__8817),
            .I(N__8812));
    InMux I__1364 (
            .O(N__8816),
            .I(N__8809));
    CascadeMux I__1363 (
            .O(N__8815),
            .I(N__8805));
    LocalMux I__1362 (
            .O(N__8812),
            .I(N__8800));
    LocalMux I__1361 (
            .O(N__8809),
            .I(N__8800));
    InMux I__1360 (
            .O(N__8808),
            .I(N__8795));
    InMux I__1359 (
            .O(N__8805),
            .I(N__8795));
    Span4Mux_h I__1358 (
            .O(N__8800),
            .I(N__8792));
    LocalMux I__1357 (
            .O(N__8795),
            .I(N__8789));
    Odrv4 I__1356 (
            .O(N__8792),
            .I(Lab_UT_rx_data_3));
    Odrv12 I__1355 (
            .O(N__8789),
            .I(Lab_UT_rx_data_3));
    CascadeMux I__1354 (
            .O(N__8784),
            .I(\Lab_UT.dictrluu0.N_103_1_cascade_ ));
    InMux I__1353 (
            .O(N__8781),
            .I(N__8778));
    LocalMux I__1352 (
            .O(N__8778),
            .I(N__8775));
    Span4Mux_h I__1351 (
            .O(N__8775),
            .I(N__8769));
    InMux I__1350 (
            .O(N__8774),
            .I(N__8766));
    InMux I__1349 (
            .O(N__8773),
            .I(N__8761));
    InMux I__1348 (
            .O(N__8772),
            .I(N__8761));
    Odrv4 I__1347 (
            .O(N__8769),
            .I(Lab_UT_rx_data_5));
    LocalMux I__1346 (
            .O(N__8766),
            .I(Lab_UT_rx_data_5));
    LocalMux I__1345 (
            .O(N__8761),
            .I(Lab_UT_rx_data_5));
    InMux I__1344 (
            .O(N__8754),
            .I(N__8751));
    LocalMux I__1343 (
            .O(N__8751),
            .I(N__8748));
    Odrv12 I__1342 (
            .O(N__8748),
            .I(\uu2.un1_w_user_lf_3Z0Z_1 ));
    CascadeMux I__1341 (
            .O(N__8745),
            .I(N__8738));
    InMux I__1340 (
            .O(N__8744),
            .I(N__8732));
    InMux I__1339 (
            .O(N__8743),
            .I(N__8732));
    InMux I__1338 (
            .O(N__8742),
            .I(N__8718));
    InMux I__1337 (
            .O(N__8741),
            .I(N__8715));
    InMux I__1336 (
            .O(N__8738),
            .I(N__8710));
    InMux I__1335 (
            .O(N__8737),
            .I(N__8710));
    LocalMux I__1334 (
            .O(N__8732),
            .I(N__8707));
    InMux I__1333 (
            .O(N__8731),
            .I(N__8700));
    InMux I__1332 (
            .O(N__8730),
            .I(N__8700));
    InMux I__1331 (
            .O(N__8729),
            .I(N__8700));
    InMux I__1330 (
            .O(N__8728),
            .I(N__8693));
    InMux I__1329 (
            .O(N__8727),
            .I(N__8693));
    InMux I__1328 (
            .O(N__8726),
            .I(N__8693));
    InMux I__1327 (
            .O(N__8725),
            .I(N__8682));
    InMux I__1326 (
            .O(N__8724),
            .I(N__8682));
    InMux I__1325 (
            .O(N__8723),
            .I(N__8682));
    InMux I__1324 (
            .O(N__8722),
            .I(N__8682));
    InMux I__1323 (
            .O(N__8721),
            .I(N__8682));
    LocalMux I__1322 (
            .O(N__8718),
            .I(Lab_UT_dspStr_cnt_1));
    LocalMux I__1321 (
            .O(N__8715),
            .I(Lab_UT_dspStr_cnt_1));
    LocalMux I__1320 (
            .O(N__8710),
            .I(Lab_UT_dspStr_cnt_1));
    Odrv12 I__1319 (
            .O(N__8707),
            .I(Lab_UT_dspStr_cnt_1));
    LocalMux I__1318 (
            .O(N__8700),
            .I(Lab_UT_dspStr_cnt_1));
    LocalMux I__1317 (
            .O(N__8693),
            .I(Lab_UT_dspStr_cnt_1));
    LocalMux I__1316 (
            .O(N__8682),
            .I(Lab_UT_dspStr_cnt_1));
    InMux I__1315 (
            .O(N__8667),
            .I(N__8661));
    CascadeMux I__1314 (
            .O(N__8666),
            .I(N__8646));
    CascadeMux I__1313 (
            .O(N__8665),
            .I(N__8643));
    InMux I__1312 (
            .O(N__8664),
            .I(N__8639));
    LocalMux I__1311 (
            .O(N__8661),
            .I(N__8636));
    InMux I__1310 (
            .O(N__8660),
            .I(N__8633));
    InMux I__1309 (
            .O(N__8659),
            .I(N__8628));
    InMux I__1308 (
            .O(N__8658),
            .I(N__8628));
    InMux I__1307 (
            .O(N__8657),
            .I(N__8625));
    InMux I__1306 (
            .O(N__8656),
            .I(N__8620));
    InMux I__1305 (
            .O(N__8655),
            .I(N__8620));
    InMux I__1304 (
            .O(N__8654),
            .I(N__8613));
    InMux I__1303 (
            .O(N__8653),
            .I(N__8613));
    InMux I__1302 (
            .O(N__8652),
            .I(N__8613));
    InMux I__1301 (
            .O(N__8651),
            .I(N__8606));
    InMux I__1300 (
            .O(N__8650),
            .I(N__8606));
    InMux I__1299 (
            .O(N__8649),
            .I(N__8606));
    InMux I__1298 (
            .O(N__8646),
            .I(N__8599));
    InMux I__1297 (
            .O(N__8643),
            .I(N__8599));
    InMux I__1296 (
            .O(N__8642),
            .I(N__8599));
    LocalMux I__1295 (
            .O(N__8639),
            .I(Lab_UT_dspStr_cnt_3));
    Odrv12 I__1294 (
            .O(N__8636),
            .I(Lab_UT_dspStr_cnt_3));
    LocalMux I__1293 (
            .O(N__8633),
            .I(Lab_UT_dspStr_cnt_3));
    LocalMux I__1292 (
            .O(N__8628),
            .I(Lab_UT_dspStr_cnt_3));
    LocalMux I__1291 (
            .O(N__8625),
            .I(Lab_UT_dspStr_cnt_3));
    LocalMux I__1290 (
            .O(N__8620),
            .I(Lab_UT_dspStr_cnt_3));
    LocalMux I__1289 (
            .O(N__8613),
            .I(Lab_UT_dspStr_cnt_3));
    LocalMux I__1288 (
            .O(N__8606),
            .I(Lab_UT_dspStr_cnt_3));
    LocalMux I__1287 (
            .O(N__8599),
            .I(Lab_UT_dspStr_cnt_3));
    CascadeMux I__1286 (
            .O(N__8580),
            .I(\uu2.mem0.N_26_1_cascade_ ));
    CascadeMux I__1285 (
            .O(N__8577),
            .I(N__8571));
    InMux I__1284 (
            .O(N__8576),
            .I(N__8555));
    InMux I__1283 (
            .O(N__8575),
            .I(N__8555));
    InMux I__1282 (
            .O(N__8574),
            .I(N__8552));
    InMux I__1281 (
            .O(N__8571),
            .I(N__8549));
    InMux I__1280 (
            .O(N__8570),
            .I(N__8546));
    InMux I__1279 (
            .O(N__8569),
            .I(N__8543));
    InMux I__1278 (
            .O(N__8568),
            .I(N__8536));
    InMux I__1277 (
            .O(N__8567),
            .I(N__8536));
    InMux I__1276 (
            .O(N__8566),
            .I(N__8536));
    InMux I__1275 (
            .O(N__8565),
            .I(N__8529));
    InMux I__1274 (
            .O(N__8564),
            .I(N__8529));
    InMux I__1273 (
            .O(N__8563),
            .I(N__8529));
    InMux I__1272 (
            .O(N__8562),
            .I(N__8522));
    InMux I__1271 (
            .O(N__8561),
            .I(N__8522));
    InMux I__1270 (
            .O(N__8560),
            .I(N__8522));
    LocalMux I__1269 (
            .O(N__8555),
            .I(N__8519));
    LocalMux I__1268 (
            .O(N__8552),
            .I(Lab_UT_dspStr_cnt_2));
    LocalMux I__1267 (
            .O(N__8549),
            .I(Lab_UT_dspStr_cnt_2));
    LocalMux I__1266 (
            .O(N__8546),
            .I(Lab_UT_dspStr_cnt_2));
    LocalMux I__1265 (
            .O(N__8543),
            .I(Lab_UT_dspStr_cnt_2));
    LocalMux I__1264 (
            .O(N__8536),
            .I(Lab_UT_dspStr_cnt_2));
    LocalMux I__1263 (
            .O(N__8529),
            .I(Lab_UT_dspStr_cnt_2));
    LocalMux I__1262 (
            .O(N__8522),
            .I(Lab_UT_dspStr_cnt_2));
    Odrv12 I__1261 (
            .O(N__8519),
            .I(Lab_UT_dspStr_cnt_2));
    CascadeMux I__1260 (
            .O(N__8502),
            .I(\resetGen.reset_count_2_i_0_a3_5Z0Z_4_cascade_ ));
    InMux I__1259 (
            .O(N__8499),
            .I(N__8496));
    LocalMux I__1258 (
            .O(N__8496),
            .I(N__8493));
    Span4Mux_v I__1257 (
            .O(N__8493),
            .I(N__8488));
    InMux I__1256 (
            .O(N__8492),
            .I(N__8483));
    InMux I__1255 (
            .O(N__8491),
            .I(N__8483));
    Odrv4 I__1254 (
            .O(N__8488),
            .I(bu_rx_data_5));
    LocalMux I__1253 (
            .O(N__8483),
            .I(bu_rx_data_5));
    InMux I__1252 (
            .O(N__8478),
            .I(N__8475));
    LocalMux I__1251 (
            .O(N__8475),
            .I(\resetGen.reset_count_2_i_0_a3_6Z0Z_4 ));
    InMux I__1250 (
            .O(N__8472),
            .I(N__8469));
    LocalMux I__1249 (
            .O(N__8469),
            .I(\resetGen.reset_count_2_i_0_a3_4Z0Z_4 ));
    InMux I__1248 (
            .O(N__8466),
            .I(N__8462));
    InMux I__1247 (
            .O(N__8465),
            .I(N__8459));
    LocalMux I__1246 (
            .O(N__8462),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    LocalMux I__1245 (
            .O(N__8459),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    CascadeMux I__1244 (
            .O(N__8454),
            .I(\buart.Z_rx.N_129_cascade_ ));
    InMux I__1243 (
            .O(N__8451),
            .I(N__8445));
    InMux I__1242 (
            .O(N__8450),
            .I(N__8445));
    LocalMux I__1241 (
            .O(N__8445),
            .I(N__8442));
    Span4Mux_v I__1240 (
            .O(N__8442),
            .I(N__8439));
    Span4Mux_h I__1239 (
            .O(N__8439),
            .I(N__8436));
    Odrv4 I__1238 (
            .O(N__8436),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    InMux I__1237 (
            .O(N__8433),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    CascadeMux I__1236 (
            .O(N__8430),
            .I(\buart.Z_rx.N_144_cascade_ ));
    InMux I__1235 (
            .O(N__8427),
            .I(N__8422));
    InMux I__1234 (
            .O(N__8426),
            .I(N__8417));
    InMux I__1233 (
            .O(N__8425),
            .I(N__8417));
    LocalMux I__1232 (
            .O(N__8422),
            .I(buart__rx_bitcount_4));
    LocalMux I__1231 (
            .O(N__8417),
            .I(buart__rx_bitcount_4));
    InMux I__1230 (
            .O(N__8412),
            .I(N__8409));
    LocalMux I__1229 (
            .O(N__8409),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    InMux I__1228 (
            .O(N__8406),
            .I(N__8400));
    InMux I__1227 (
            .O(N__8405),
            .I(N__8397));
    InMux I__1226 (
            .O(N__8404),
            .I(N__8392));
    InMux I__1225 (
            .O(N__8403),
            .I(N__8392));
    LocalMux I__1224 (
            .O(N__8400),
            .I(buart__rx_bitcount_1));
    LocalMux I__1223 (
            .O(N__8397),
            .I(buart__rx_bitcount_1));
    LocalMux I__1222 (
            .O(N__8392),
            .I(buart__rx_bitcount_1));
    CascadeMux I__1221 (
            .O(N__8385),
            .I(N__8382));
    InMux I__1220 (
            .O(N__8382),
            .I(N__8379));
    LocalMux I__1219 (
            .O(N__8379),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__1218 (
            .O(N__8376),
            .I(N__8373));
    LocalMux I__1217 (
            .O(N__8373),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    IoInMux I__1216 (
            .O(N__8370),
            .I(N__8366));
    CascadeMux I__1215 (
            .O(N__8369),
            .I(N__8363));
    LocalMux I__1214 (
            .O(N__8366),
            .I(N__8360));
    InMux I__1213 (
            .O(N__8363),
            .I(N__8357));
    Span4Mux_s1_v I__1212 (
            .O(N__8360),
            .I(N__8354));
    LocalMux I__1211 (
            .O(N__8357),
            .I(N__8351));
    Odrv4 I__1210 (
            .O(N__8354),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__1209 (
            .O(N__8351),
            .I(CONSTANT_ONE_NET));
    InMux I__1208 (
            .O(N__8346),
            .I(N__8343));
    LocalMux I__1207 (
            .O(N__8343),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__1206 (
            .O(N__8340),
            .I(N__8337));
    LocalMux I__1205 (
            .O(N__8337),
            .I(N__8334));
    Span4Mux_v I__1204 (
            .O(N__8334),
            .I(N__8331));
    Odrv4 I__1203 (
            .O(N__8331),
            .I(vbuf_tx_data_3));
    InMux I__1202 (
            .O(N__8328),
            .I(N__8325));
    LocalMux I__1201 (
            .O(N__8325),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__1200 (
            .O(N__8322),
            .I(N__8319));
    LocalMux I__1199 (
            .O(N__8319),
            .I(vbuf_tx_data_4));
    InMux I__1198 (
            .O(N__8316),
            .I(N__8313));
    LocalMux I__1197 (
            .O(N__8313),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__1196 (
            .O(N__8310),
            .I(N__8307));
    LocalMux I__1195 (
            .O(N__8307),
            .I(vbuf_tx_data_5));
    InMux I__1194 (
            .O(N__8304),
            .I(N__8301));
    LocalMux I__1193 (
            .O(N__8301),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    InMux I__1192 (
            .O(N__8298),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__1191 (
            .O(N__8295),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    InMux I__1190 (
            .O(N__8292),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__1189 (
            .O(N__8289),
            .I(N__8286));
    LocalMux I__1188 (
            .O(N__8286),
            .I(N__8283));
    Odrv4 I__1187 (
            .O(N__8283),
            .I(\uu2.r_data_wire_4 ));
    InMux I__1186 (
            .O(N__8280),
            .I(N__8277));
    LocalMux I__1185 (
            .O(N__8277),
            .I(N__8274));
    Odrv4 I__1184 (
            .O(N__8274),
            .I(\uu2.r_data_wire_5 ));
    InMux I__1183 (
            .O(N__8271),
            .I(N__8268));
    LocalMux I__1182 (
            .O(N__8268),
            .I(N__8265));
    Odrv4 I__1181 (
            .O(N__8265),
            .I(\uu2.r_data_wire_6 ));
    InMux I__1180 (
            .O(N__8262),
            .I(N__8259));
    LocalMux I__1179 (
            .O(N__8259),
            .I(N__8256));
    Odrv4 I__1178 (
            .O(N__8256),
            .I(\uu2.r_data_wire_7 ));
    CascadeMux I__1177 (
            .O(N__8253),
            .I(N__8250));
    InMux I__1176 (
            .O(N__8250),
            .I(N__8247));
    LocalMux I__1175 (
            .O(N__8247),
            .I(vbuf_tx_data_0));
    InMux I__1174 (
            .O(N__8244),
            .I(N__8241));
    LocalMux I__1173 (
            .O(N__8241),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__1172 (
            .O(N__8238),
            .I(N__8235));
    LocalMux I__1171 (
            .O(N__8235),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__1170 (
            .O(N__8232),
            .I(N__8229));
    LocalMux I__1169 (
            .O(N__8229),
            .I(N__8226));
    Span4Mux_s3_h I__1168 (
            .O(N__8226),
            .I(N__8223));
    Odrv4 I__1167 (
            .O(N__8223),
            .I(o_serial_data_c));
    InMux I__1166 (
            .O(N__8220),
            .I(N__8217));
    LocalMux I__1165 (
            .O(N__8217),
            .I(vbuf_tx_data_1));
    InMux I__1164 (
            .O(N__8214),
            .I(N__8211));
    LocalMux I__1163 (
            .O(N__8211),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__1162 (
            .O(N__8208),
            .I(N__8205));
    LocalMux I__1161 (
            .O(N__8205),
            .I(vbuf_tx_data_2));
    InMux I__1160 (
            .O(N__8202),
            .I(N__8199));
    LocalMux I__1159 (
            .O(N__8199),
            .I(\uu2.bitmap_pmux_1_1_a8_1_2_0 ));
    InMux I__1158 (
            .O(N__8196),
            .I(N__8193));
    LocalMux I__1157 (
            .O(N__8193),
            .I(\uu2.N_326_0 ));
    CascadeMux I__1156 (
            .O(N__8190),
            .I(\uu2.bitmap_pmux_1_1_a8_1_1_cascade_ ));
    InMux I__1155 (
            .O(N__8187),
            .I(N__8184));
    LocalMux I__1154 (
            .O(N__8184),
            .I(\uu2.bitmap_pmux_1_1_a8_0_1 ));
    InMux I__1153 (
            .O(N__8181),
            .I(N__8178));
    LocalMux I__1152 (
            .O(N__8178),
            .I(\uu2.bitmap_pmux_1_1_1_tz ));
    CascadeMux I__1151 (
            .O(N__8175),
            .I(\uu2.bitmap_pmux_1_1_1_tz_cascade_ ));
    CascadeMux I__1150 (
            .O(N__8172),
            .I(N__8169));
    InMux I__1149 (
            .O(N__8169),
            .I(N__8166));
    LocalMux I__1148 (
            .O(N__8166),
            .I(N__8163));
    Span4Mux_v I__1147 (
            .O(N__8163),
            .I(N__8159));
    InMux I__1146 (
            .O(N__8162),
            .I(N__8156));
    Odrv4 I__1145 (
            .O(N__8159),
            .I(L3_tx_data_3));
    LocalMux I__1144 (
            .O(N__8156),
            .I(L3_tx_data_3));
    InMux I__1143 (
            .O(N__8151),
            .I(N__8148));
    LocalMux I__1142 (
            .O(N__8148),
            .I(N__8145));
    Odrv4 I__1141 (
            .O(N__8145),
            .I(\uu2.mem0.w_data_1_0_0_3 ));
    IoInMux I__1140 (
            .O(N__8142),
            .I(N__8138));
    InMux I__1139 (
            .O(N__8141),
            .I(N__8135));
    LocalMux I__1138 (
            .O(N__8138),
            .I(N__8132));
    LocalMux I__1137 (
            .O(N__8135),
            .I(N__8129));
    Span12Mux_s5_v I__1136 (
            .O(N__8132),
            .I(N__8124));
    Span12Mux_s5_h I__1135 (
            .O(N__8129),
            .I(N__8124));
    Odrv12 I__1134 (
            .O(N__8124),
            .I(latticehx1k_pll_inst_PLLOUTCORE_i));
    CEMux I__1133 (
            .O(N__8121),
            .I(N__8117));
    SRMux I__1132 (
            .O(N__8120),
            .I(N__8114));
    LocalMux I__1131 (
            .O(N__8117),
            .I(N__8111));
    LocalMux I__1130 (
            .O(N__8114),
            .I(N__8108));
    Span4Mux_v I__1129 (
            .O(N__8111),
            .I(N__8105));
    Odrv4 I__1128 (
            .O(N__8108),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    Odrv4 I__1127 (
            .O(N__8105),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    InMux I__1126 (
            .O(N__8100),
            .I(N__8097));
    LocalMux I__1125 (
            .O(N__8097),
            .I(N__8090));
    CascadeMux I__1124 (
            .O(N__8096),
            .I(N__8087));
    CascadeMux I__1123 (
            .O(N__8095),
            .I(N__8084));
    InMux I__1122 (
            .O(N__8094),
            .I(N__8077));
    InMux I__1121 (
            .O(N__8093),
            .I(N__8077));
    Span4Mux_v I__1120 (
            .O(N__8090),
            .I(N__8074));
    InMux I__1119 (
            .O(N__8087),
            .I(N__8065));
    InMux I__1118 (
            .O(N__8084),
            .I(N__8065));
    InMux I__1117 (
            .O(N__8083),
            .I(N__8065));
    InMux I__1116 (
            .O(N__8082),
            .I(N__8065));
    LocalMux I__1115 (
            .O(N__8077),
            .I(\uu2.w_addr_userZ0Z_0 ));
    Odrv4 I__1114 (
            .O(N__8074),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__1113 (
            .O(N__8065),
            .I(\uu2.w_addr_userZ0Z_0 ));
    CascadeMux I__1112 (
            .O(N__8058),
            .I(N__8055));
    InMux I__1111 (
            .O(N__8055),
            .I(N__8052));
    LocalMux I__1110 (
            .O(N__8052),
            .I(N__8049));
    Odrv4 I__1109 (
            .O(N__8049),
            .I(\uu2.mem0.w_addr_0 ));
    InMux I__1108 (
            .O(N__8046),
            .I(N__8043));
    LocalMux I__1107 (
            .O(N__8043),
            .I(N__8040));
    Odrv4 I__1106 (
            .O(N__8040),
            .I(\uu2.r_data_wire_1 ));
    InMux I__1105 (
            .O(N__8037),
            .I(N__8034));
    LocalMux I__1104 (
            .O(N__8034),
            .I(N__8031));
    Odrv4 I__1103 (
            .O(N__8031),
            .I(\uu2.r_data_wire_2 ));
    InMux I__1102 (
            .O(N__8028),
            .I(N__8025));
    LocalMux I__1101 (
            .O(N__8025),
            .I(N__8022));
    Span4Mux_v I__1100 (
            .O(N__8022),
            .I(N__8019));
    Odrv4 I__1099 (
            .O(N__8019),
            .I(\uu2.r_data_wire_0 ));
    CascadeMux I__1098 (
            .O(N__8016),
            .I(\uu2.mem0.N_7_0_cascade_ ));
    InMux I__1097 (
            .O(N__8013),
            .I(N__8010));
    LocalMux I__1096 (
            .O(N__8010),
            .I(\uu2.mem0.w_data_1 ));
    InMux I__1095 (
            .O(N__8007),
            .I(N__8004));
    LocalMux I__1094 (
            .O(N__8004),
            .I(N__8001));
    Odrv4 I__1093 (
            .O(N__8001),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_22 ));
    CascadeMux I__1092 (
            .O(N__7998),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_ ));
    InMux I__1091 (
            .O(N__7995),
            .I(N__7992));
    LocalMux I__1090 (
            .O(N__7992),
            .I(\uu2.mem0.w_data_4 ));
    CascadeMux I__1089 (
            .O(N__7989),
            .I(N__7986));
    InMux I__1088 (
            .O(N__7986),
            .I(N__7983));
    LocalMux I__1087 (
            .O(N__7983),
            .I(\uu2.mem0.G_14_0_a6_0_0_1 ));
    InMux I__1086 (
            .O(N__7980),
            .I(N__7977));
    LocalMux I__1085 (
            .O(N__7977),
            .I(\uu2.mem0.w_data_3 ));
    CascadeMux I__1084 (
            .O(N__7974),
            .I(\uu2.N_326_0_cascade_ ));
    CascadeMux I__1083 (
            .O(N__7971),
            .I(\uu2.vbuf_raddr.un469_ci_0_cascade_ ));
    CascadeMux I__1082 (
            .O(N__7968),
            .I(N__7965));
    InMux I__1081 (
            .O(N__7965),
            .I(N__7962));
    LocalMux I__1080 (
            .O(N__7962),
            .I(N__7958));
    InMux I__1079 (
            .O(N__7961),
            .I(N__7955));
    Odrv4 I__1078 (
            .O(N__7958),
            .I(\uu2.r_addrZ0Z_8 ));
    LocalMux I__1077 (
            .O(N__7955),
            .I(\uu2.r_addrZ0Z_8 ));
    CascadeMux I__1076 (
            .O(N__7950),
            .I(N__7947));
    InMux I__1075 (
            .O(N__7947),
            .I(N__7944));
    LocalMux I__1074 (
            .O(N__7944),
            .I(N__7941));
    Span4Mux_h I__1073 (
            .O(N__7941),
            .I(N__7935));
    InMux I__1072 (
            .O(N__7940),
            .I(N__7932));
    InMux I__1071 (
            .O(N__7939),
            .I(N__7927));
    InMux I__1070 (
            .O(N__7938),
            .I(N__7927));
    Odrv4 I__1069 (
            .O(N__7935),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__1068 (
            .O(N__7932),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__1067 (
            .O(N__7927),
            .I(\uu2.r_addrZ0Z_5 ));
    CascadeMux I__1066 (
            .O(N__7920),
            .I(N__7915));
    CascadeMux I__1065 (
            .O(N__7919),
            .I(N__7911));
    InMux I__1064 (
            .O(N__7918),
            .I(N__7908));
    InMux I__1063 (
            .O(N__7915),
            .I(N__7905));
    InMux I__1062 (
            .O(N__7914),
            .I(N__7899));
    InMux I__1061 (
            .O(N__7911),
            .I(N__7899));
    LocalMux I__1060 (
            .O(N__7908),
            .I(N__7894));
    LocalMux I__1059 (
            .O(N__7905),
            .I(N__7894));
    InMux I__1058 (
            .O(N__7904),
            .I(N__7891));
    LocalMux I__1057 (
            .O(N__7899),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__1056 (
            .O(N__7894),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__1055 (
            .O(N__7891),
            .I(\uu2.r_addrZ0Z_4 ));
    InMux I__1054 (
            .O(N__7884),
            .I(N__7881));
    LocalMux I__1053 (
            .O(N__7881),
            .I(\uu2.vbuf_raddr.un447_ci_3 ));
    CascadeMux I__1052 (
            .O(N__7878),
            .I(N__7875));
    InMux I__1051 (
            .O(N__7875),
            .I(N__7872));
    LocalMux I__1050 (
            .O(N__7872),
            .I(N__7866));
    InMux I__1049 (
            .O(N__7871),
            .I(N__7863));
    InMux I__1048 (
            .O(N__7870),
            .I(N__7858));
    InMux I__1047 (
            .O(N__7869),
            .I(N__7858));
    Odrv4 I__1046 (
            .O(N__7866),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1045 (
            .O(N__7863),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1044 (
            .O(N__7858),
            .I(\uu2.r_addrZ0Z_6 ));
    CascadeMux I__1043 (
            .O(N__7851),
            .I(\uu2.vbuf_raddr.un447_ci_3_cascade_ ));
    InMux I__1042 (
            .O(N__7848),
            .I(N__7840));
    InMux I__1041 (
            .O(N__7847),
            .I(N__7840));
    InMux I__1040 (
            .O(N__7846),
            .I(N__7835));
    InMux I__1039 (
            .O(N__7845),
            .I(N__7835));
    LocalMux I__1038 (
            .O(N__7840),
            .I(\uu2.un425_ci_0 ));
    LocalMux I__1037 (
            .O(N__7835),
            .I(\uu2.un425_ci_0 ));
    CascadeMux I__1036 (
            .O(N__7830),
            .I(N__7827));
    InMux I__1035 (
            .O(N__7827),
            .I(N__7824));
    LocalMux I__1034 (
            .O(N__7824),
            .I(N__7819));
    InMux I__1033 (
            .O(N__7823),
            .I(N__7816));
    InMux I__1032 (
            .O(N__7822),
            .I(N__7813));
    Odrv4 I__1031 (
            .O(N__7819),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__1030 (
            .O(N__7816),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__1029 (
            .O(N__7813),
            .I(\uu2.r_addrZ0Z_7 ));
    CascadeMux I__1028 (
            .O(N__7806),
            .I(N__7803));
    InMux I__1027 (
            .O(N__7803),
            .I(N__7798));
    CascadeMux I__1026 (
            .O(N__7802),
            .I(N__7795));
    CascadeMux I__1025 (
            .O(N__7801),
            .I(N__7792));
    LocalMux I__1024 (
            .O(N__7798),
            .I(N__7789));
    InMux I__1023 (
            .O(N__7795),
            .I(N__7784));
    InMux I__1022 (
            .O(N__7792),
            .I(N__7784));
    Odrv4 I__1021 (
            .O(N__7789),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__1020 (
            .O(N__7784),
            .I(\uu2.r_addrZ0Z_3 ));
    InMux I__1019 (
            .O(N__7779),
            .I(N__7776));
    LocalMux I__1018 (
            .O(N__7776),
            .I(N__7773));
    Odrv4 I__1017 (
            .O(N__7773),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_21 ));
    InMux I__1016 (
            .O(N__7770),
            .I(N__7767));
    LocalMux I__1015 (
            .O(N__7767),
            .I(\uu2.mem0.w_data_0 ));
    InMux I__1014 (
            .O(N__7764),
            .I(N__7761));
    LocalMux I__1013 (
            .O(N__7761),
            .I(N__7758));
    Span4Mux_v I__1012 (
            .O(N__7758),
            .I(N__7755));
    Odrv4 I__1011 (
            .O(N__7755),
            .I(\uu2.mem0.w_data_ns_1_5 ));
    InMux I__1010 (
            .O(N__7752),
            .I(N__7749));
    LocalMux I__1009 (
            .O(N__7749),
            .I(\uu2.mem0.w_data_5 ));
    InMux I__1008 (
            .O(N__7746),
            .I(N__7743));
    LocalMux I__1007 (
            .O(N__7743),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_17 ));
    CascadeMux I__1006 (
            .O(N__7740),
            .I(\uu2.mem0.G_14_0_a6_0_cascade_ ));
    CascadeMux I__1005 (
            .O(N__7737),
            .I(N__7734));
    InMux I__1004 (
            .O(N__7734),
            .I(N__7730));
    InMux I__1003 (
            .O(N__7733),
            .I(N__7727));
    LocalMux I__1002 (
            .O(N__7730),
            .I(N__7721));
    LocalMux I__1001 (
            .O(N__7727),
            .I(N__7721));
    InMux I__1000 (
            .O(N__7726),
            .I(N__7717));
    Span4Mux_v I__999 (
            .O(N__7721),
            .I(N__7714));
    InMux I__998 (
            .O(N__7720),
            .I(N__7711));
    LocalMux I__997 (
            .O(N__7717),
            .I(\Lab_UT.secuu0.un197_ci_9 ));
    Odrv4 I__996 (
            .O(N__7714),
            .I(\Lab_UT.secuu0.un197_ci_9 ));
    LocalMux I__995 (
            .O(N__7711),
            .I(\Lab_UT.secuu0.un197_ci_9 ));
    InMux I__994 (
            .O(N__7704),
            .I(N__7699));
    InMux I__993 (
            .O(N__7703),
            .I(N__7696));
    InMux I__992 (
            .O(N__7702),
            .I(N__7693));
    LocalMux I__991 (
            .O(N__7699),
            .I(N__7690));
    LocalMux I__990 (
            .O(N__7696),
            .I(\Lab_UT.secuu0.l_countZ0Z_12 ));
    LocalMux I__989 (
            .O(N__7693),
            .I(\Lab_UT.secuu0.l_countZ0Z_12 ));
    Odrv4 I__988 (
            .O(N__7690),
            .I(\Lab_UT.secuu0.l_countZ0Z_12 ));
    InMux I__987 (
            .O(N__7683),
            .I(N__7677));
    InMux I__986 (
            .O(N__7682),
            .I(N__7677));
    LocalMux I__985 (
            .O(N__7677),
            .I(N__7667));
    InMux I__984 (
            .O(N__7676),
            .I(N__7662));
    InMux I__983 (
            .O(N__7675),
            .I(N__7662));
    InMux I__982 (
            .O(N__7674),
            .I(N__7659));
    InMux I__981 (
            .O(N__7673),
            .I(N__7654));
    InMux I__980 (
            .O(N__7672),
            .I(N__7654));
    InMux I__979 (
            .O(N__7671),
            .I(N__7650));
    CascadeMux I__978 (
            .O(N__7670),
            .I(N__7647));
    Span4Mux_v I__977 (
            .O(N__7667),
            .I(N__7637));
    LocalMux I__976 (
            .O(N__7662),
            .I(N__7637));
    LocalMux I__975 (
            .O(N__7659),
            .I(N__7637));
    LocalMux I__974 (
            .O(N__7654),
            .I(N__7637));
    InMux I__973 (
            .O(N__7653),
            .I(N__7634));
    LocalMux I__972 (
            .O(N__7650),
            .I(N__7631));
    InMux I__971 (
            .O(N__7647),
            .I(N__7626));
    InMux I__970 (
            .O(N__7646),
            .I(N__7626));
    Span4Mux_h I__969 (
            .O(N__7637),
            .I(N__7623));
    LocalMux I__968 (
            .O(N__7634),
            .I(N__7620));
    Odrv4 I__967 (
            .O(N__7631),
            .I(\Lab_UT.secuu0.un153_ci ));
    LocalMux I__966 (
            .O(N__7626),
            .I(\Lab_UT.secuu0.un153_ci ));
    Odrv4 I__965 (
            .O(N__7623),
            .I(\Lab_UT.secuu0.un153_ci ));
    Odrv12 I__964 (
            .O(N__7620),
            .I(\Lab_UT.secuu0.un153_ci ));
    InMux I__963 (
            .O(N__7611),
            .I(N__7608));
    LocalMux I__962 (
            .O(N__7608),
            .I(\Lab_UT.secuu0.un208_ci_0 ));
    CascadeMux I__961 (
            .O(N__7605),
            .I(N__7601));
    InMux I__960 (
            .O(N__7604),
            .I(N__7598));
    InMux I__959 (
            .O(N__7601),
            .I(N__7595));
    LocalMux I__958 (
            .O(N__7598),
            .I(N__7592));
    LocalMux I__957 (
            .O(N__7595),
            .I(\Lab_UT.secuu0.l_countZ0Z_13 ));
    Odrv4 I__956 (
            .O(N__7592),
            .I(\Lab_UT.secuu0.l_countZ0Z_13 ));
    CEMux I__955 (
            .O(N__7587),
            .I(N__7566));
    CEMux I__954 (
            .O(N__7586),
            .I(N__7566));
    CEMux I__953 (
            .O(N__7585),
            .I(N__7566));
    CEMux I__952 (
            .O(N__7584),
            .I(N__7566));
    CEMux I__951 (
            .O(N__7583),
            .I(N__7566));
    CEMux I__950 (
            .O(N__7582),
            .I(N__7566));
    CEMux I__949 (
            .O(N__7581),
            .I(N__7566));
    GlobalMux I__948 (
            .O(N__7566),
            .I(N__7563));
    gio2CtrlBuf I__947 (
            .O(N__7563),
            .I(\Lab_UT.secuu0.un11_l_count_i_g ));
    CascadeMux I__946 (
            .O(N__7560),
            .I(N__7557));
    InMux I__945 (
            .O(N__7557),
            .I(N__7546));
    InMux I__944 (
            .O(N__7556),
            .I(N__7546));
    InMux I__943 (
            .O(N__7555),
            .I(N__7546));
    InMux I__942 (
            .O(N__7554),
            .I(N__7541));
    InMux I__941 (
            .O(N__7553),
            .I(N__7541));
    LocalMux I__940 (
            .O(N__7546),
            .I(N__7535));
    LocalMux I__939 (
            .O(N__7541),
            .I(N__7535));
    InMux I__938 (
            .O(N__7540),
            .I(N__7532));
    Span4Mux_h I__937 (
            .O(N__7535),
            .I(N__7529));
    LocalMux I__936 (
            .O(N__7532),
            .I(\Lab_UT.secuu0.l_precountZ0Z_0 ));
    Odrv4 I__935 (
            .O(N__7529),
            .I(\Lab_UT.secuu0.l_precountZ0Z_0 ));
    CascadeMux I__934 (
            .O(N__7524),
            .I(\uu2.un425_ci_0_cascade_ ));
    InMux I__933 (
            .O(N__7521),
            .I(N__7518));
    LocalMux I__932 (
            .O(N__7518),
            .I(N__7512));
    InMux I__931 (
            .O(N__7517),
            .I(N__7507));
    InMux I__930 (
            .O(N__7516),
            .I(N__7507));
    InMux I__929 (
            .O(N__7515),
            .I(N__7504));
    Odrv4 I__928 (
            .O(N__7512),
            .I(\Lab_UT.secuu0.l_countZ0Z_10 ));
    LocalMux I__927 (
            .O(N__7507),
            .I(\Lab_UT.secuu0.l_countZ0Z_10 ));
    LocalMux I__926 (
            .O(N__7504),
            .I(\Lab_UT.secuu0.l_countZ0Z_10 ));
    CascadeMux I__925 (
            .O(N__7497),
            .I(\Lab_UT.secuu0.un186_ci_0_cascade_ ));
    InMux I__924 (
            .O(N__7494),
            .I(N__7490));
    InMux I__923 (
            .O(N__7493),
            .I(N__7485));
    LocalMux I__922 (
            .O(N__7490),
            .I(N__7480));
    InMux I__921 (
            .O(N__7489),
            .I(N__7477));
    InMux I__920 (
            .O(N__7488),
            .I(N__7474));
    LocalMux I__919 (
            .O(N__7485),
            .I(N__7471));
    InMux I__918 (
            .O(N__7484),
            .I(N__7466));
    InMux I__917 (
            .O(N__7483),
            .I(N__7466));
    Span4Mux_s3_v I__916 (
            .O(N__7480),
            .I(N__7457));
    LocalMux I__915 (
            .O(N__7477),
            .I(N__7457));
    LocalMux I__914 (
            .O(N__7474),
            .I(N__7457));
    Span4Mux_v I__913 (
            .O(N__7471),
            .I(N__7457));
    LocalMux I__912 (
            .O(N__7466),
            .I(\Lab_UT.secuu0.l_countZ0Z_8 ));
    Odrv4 I__911 (
            .O(N__7457),
            .I(\Lab_UT.secuu0.l_countZ0Z_8 ));
    InMux I__910 (
            .O(N__7452),
            .I(N__7448));
    InMux I__909 (
            .O(N__7451),
            .I(N__7445));
    LocalMux I__908 (
            .O(N__7448),
            .I(N__7441));
    LocalMux I__907 (
            .O(N__7445),
            .I(N__7436));
    InMux I__906 (
            .O(N__7444),
            .I(N__7433));
    Span4Mux_h I__905 (
            .O(N__7441),
            .I(N__7430));
    InMux I__904 (
            .O(N__7440),
            .I(N__7425));
    InMux I__903 (
            .O(N__7439),
            .I(N__7425));
    Span4Mux_h I__902 (
            .O(N__7436),
            .I(N__7422));
    LocalMux I__901 (
            .O(N__7433),
            .I(\Lab_UT.secuu0.l_countZ0Z_9 ));
    Odrv4 I__900 (
            .O(N__7430),
            .I(\Lab_UT.secuu0.l_countZ0Z_9 ));
    LocalMux I__899 (
            .O(N__7425),
            .I(\Lab_UT.secuu0.l_countZ0Z_9 ));
    Odrv4 I__898 (
            .O(N__7422),
            .I(\Lab_UT.secuu0.l_countZ0Z_9 ));
    InMux I__897 (
            .O(N__7413),
            .I(N__7408));
    InMux I__896 (
            .O(N__7412),
            .I(N__7403));
    InMux I__895 (
            .O(N__7411),
            .I(N__7403));
    LocalMux I__894 (
            .O(N__7408),
            .I(N__7400));
    LocalMux I__893 (
            .O(N__7403),
            .I(\Lab_UT.secuu0.l_countZ0Z_7 ));
    Odrv4 I__892 (
            .O(N__7400),
            .I(\Lab_UT.secuu0.l_countZ0Z_7 ));
    CascadeMux I__891 (
            .O(N__7395),
            .I(N__7391));
    InMux I__890 (
            .O(N__7394),
            .I(N__7387));
    InMux I__889 (
            .O(N__7391),
            .I(N__7384));
    InMux I__888 (
            .O(N__7390),
            .I(N__7381));
    LocalMux I__887 (
            .O(N__7387),
            .I(N__7378));
    LocalMux I__886 (
            .O(N__7384),
            .I(\Lab_UT.secuu0.l_countZ0Z_3 ));
    LocalMux I__885 (
            .O(N__7381),
            .I(\Lab_UT.secuu0.l_countZ0Z_3 ));
    Odrv4 I__884 (
            .O(N__7378),
            .I(\Lab_UT.secuu0.l_countZ0Z_3 ));
    CascadeMux I__883 (
            .O(N__7371),
            .I(N__7368));
    InMux I__882 (
            .O(N__7368),
            .I(N__7364));
    InMux I__881 (
            .O(N__7367),
            .I(N__7360));
    LocalMux I__880 (
            .O(N__7364),
            .I(N__7357));
    InMux I__879 (
            .O(N__7363),
            .I(N__7354));
    LocalMux I__878 (
            .O(N__7360),
            .I(\Lab_UT.secuu0.l_countZ0Z_11 ));
    Odrv4 I__877 (
            .O(N__7357),
            .I(\Lab_UT.secuu0.l_countZ0Z_11 ));
    LocalMux I__876 (
            .O(N__7354),
            .I(\Lab_UT.secuu0.l_countZ0Z_11 ));
    CascadeMux I__875 (
            .O(N__7347),
            .I(\Lab_UT.secuu0.un4_l_count_11_cascade_ ));
    InMux I__874 (
            .O(N__7344),
            .I(N__7338));
    InMux I__873 (
            .O(N__7343),
            .I(N__7335));
    InMux I__872 (
            .O(N__7342),
            .I(N__7330));
    InMux I__871 (
            .O(N__7341),
            .I(N__7330));
    LocalMux I__870 (
            .O(N__7338),
            .I(N__7327));
    LocalMux I__869 (
            .O(N__7335),
            .I(\Lab_UT.secuu0.l_countZ0Z_6 ));
    LocalMux I__868 (
            .O(N__7330),
            .I(\Lab_UT.secuu0.l_countZ0Z_6 ));
    Odrv4 I__867 (
            .O(N__7327),
            .I(\Lab_UT.secuu0.l_countZ0Z_6 ));
    InMux I__866 (
            .O(N__7320),
            .I(N__7317));
    LocalMux I__865 (
            .O(N__7317),
            .I(N__7314));
    Odrv4 I__864 (
            .O(N__7314),
            .I(\Lab_UT.secuu0.un4_l_count_16 ));
    CascadeMux I__863 (
            .O(N__7311),
            .I(N__7307));
    CascadeMux I__862 (
            .O(N__7310),
            .I(N__7303));
    InMux I__861 (
            .O(N__7307),
            .I(N__7300));
    InMux I__860 (
            .O(N__7306),
            .I(N__7295));
    InMux I__859 (
            .O(N__7303),
            .I(N__7295));
    LocalMux I__858 (
            .O(N__7300),
            .I(\Lab_UT.secuu0.l_countZ0Z_17 ));
    LocalMux I__857 (
            .O(N__7295),
            .I(\Lab_UT.secuu0.l_countZ0Z_17 ));
    CascadeMux I__856 (
            .O(N__7290),
            .I(N__7285));
    InMux I__855 (
            .O(N__7289),
            .I(N__7282));
    InMux I__854 (
            .O(N__7288),
            .I(N__7277));
    InMux I__853 (
            .O(N__7285),
            .I(N__7277));
    LocalMux I__852 (
            .O(N__7282),
            .I(N__7274));
    LocalMux I__851 (
            .O(N__7277),
            .I(N__7271));
    Span4Mux_h I__850 (
            .O(N__7274),
            .I(N__7268));
    Odrv4 I__849 (
            .O(N__7271),
            .I(\Lab_UT.secuu0.un241_ci_2 ));
    Odrv4 I__848 (
            .O(N__7268),
            .I(\Lab_UT.secuu0.un241_ci_2 ));
    InMux I__847 (
            .O(N__7263),
            .I(N__7259));
    CascadeMux I__846 (
            .O(N__7262),
            .I(N__7254));
    LocalMux I__845 (
            .O(N__7259),
            .I(N__7251));
    InMux I__844 (
            .O(N__7258),
            .I(N__7246));
    InMux I__843 (
            .O(N__7257),
            .I(N__7246));
    InMux I__842 (
            .O(N__7254),
            .I(N__7243));
    Span4Mux_v I__841 (
            .O(N__7251),
            .I(N__7240));
    LocalMux I__840 (
            .O(N__7246),
            .I(\Lab_UT.secuu0.l_countZ0Z_16 ));
    LocalMux I__839 (
            .O(N__7243),
            .I(\Lab_UT.secuu0.l_countZ0Z_16 ));
    Odrv4 I__838 (
            .O(N__7240),
            .I(\Lab_UT.secuu0.l_countZ0Z_16 ));
    InMux I__837 (
            .O(N__7233),
            .I(N__7230));
    LocalMux I__836 (
            .O(N__7230),
            .I(\Lab_UT.secuu0.un263_ci ));
    InMux I__835 (
            .O(N__7227),
            .I(N__7223));
    InMux I__834 (
            .O(N__7226),
            .I(N__7220));
    LocalMux I__833 (
            .O(N__7223),
            .I(\Lab_UT.secuu0.l_countZ0Z_18 ));
    LocalMux I__832 (
            .O(N__7220),
            .I(\Lab_UT.secuu0.l_countZ0Z_18 ));
    CascadeMux I__831 (
            .O(N__7215),
            .I(\uu2.un2_w_addr_user_5_cascade_ ));
    InMux I__830 (
            .O(N__7212),
            .I(N__7209));
    LocalMux I__829 (
            .O(N__7209),
            .I(\uu2.un2_w_addr_user_4 ));
    InMux I__828 (
            .O(N__7206),
            .I(N__7203));
    LocalMux I__827 (
            .O(N__7203),
            .I(N__7200));
    Odrv4 I__826 (
            .O(N__7200),
            .I(\uu2.un2_w_addr_user ));
    InMux I__825 (
            .O(N__7197),
            .I(N__7180));
    InMux I__824 (
            .O(N__7196),
            .I(N__7180));
    InMux I__823 (
            .O(N__7195),
            .I(N__7180));
    InMux I__822 (
            .O(N__7194),
            .I(N__7180));
    InMux I__821 (
            .O(N__7193),
            .I(N__7169));
    InMux I__820 (
            .O(N__7192),
            .I(N__7169));
    InMux I__819 (
            .O(N__7191),
            .I(N__7169));
    InMux I__818 (
            .O(N__7190),
            .I(N__7169));
    InMux I__817 (
            .O(N__7189),
            .I(N__7169));
    LocalMux I__816 (
            .O(N__7180),
            .I(\uu2.un27_w_addr_user_i ));
    LocalMux I__815 (
            .O(N__7169),
            .I(\uu2.un27_w_addr_user_i ));
    SRMux I__814 (
            .O(N__7164),
            .I(N__7161));
    LocalMux I__813 (
            .O(N__7161),
            .I(N__7157));
    SRMux I__812 (
            .O(N__7160),
            .I(N__7154));
    Span4Mux_v I__811 (
            .O(N__7157),
            .I(N__7151));
    LocalMux I__810 (
            .O(N__7154),
            .I(N__7148));
    Odrv4 I__809 (
            .O(N__7151),
            .I(\uu2.w_addr_user_RNIKHHELZ0Z_2 ));
    Odrv4 I__808 (
            .O(N__7148),
            .I(\uu2.w_addr_user_RNIKHHELZ0Z_2 ));
    CascadeMux I__807 (
            .O(N__7143),
            .I(N__7140));
    InMux I__806 (
            .O(N__7140),
            .I(N__7137));
    LocalMux I__805 (
            .O(N__7137),
            .I(\uu2.o_adder_vbuf_w_addr_user_3 ));
    InMux I__804 (
            .O(N__7134),
            .I(N__7124));
    InMux I__803 (
            .O(N__7133),
            .I(N__7124));
    InMux I__802 (
            .O(N__7132),
            .I(N__7121));
    InMux I__801 (
            .O(N__7131),
            .I(N__7118));
    InMux I__800 (
            .O(N__7130),
            .I(N__7115));
    InMux I__799 (
            .O(N__7129),
            .I(N__7112));
    LocalMux I__798 (
            .O(N__7124),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__797 (
            .O(N__7121),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__796 (
            .O(N__7118),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__795 (
            .O(N__7115),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__794 (
            .O(N__7112),
            .I(\uu2.w_addr_userZ0Z_1 ));
    CascadeMux I__793 (
            .O(N__7101),
            .I(N__7096));
    InMux I__792 (
            .O(N__7100),
            .I(N__7089));
    InMux I__791 (
            .O(N__7099),
            .I(N__7089));
    InMux I__790 (
            .O(N__7096),
            .I(N__7086));
    InMux I__789 (
            .O(N__7095),
            .I(N__7083));
    InMux I__788 (
            .O(N__7094),
            .I(N__7080));
    LocalMux I__787 (
            .O(N__7089),
            .I(\uu2.un425_ci ));
    LocalMux I__786 (
            .O(N__7086),
            .I(\uu2.un425_ci ));
    LocalMux I__785 (
            .O(N__7083),
            .I(\uu2.un425_ci ));
    LocalMux I__784 (
            .O(N__7080),
            .I(\uu2.un425_ci ));
    InMux I__783 (
            .O(N__7071),
            .I(N__7068));
    LocalMux I__782 (
            .O(N__7068),
            .I(N__7065));
    Odrv4 I__781 (
            .O(N__7065),
            .I(\uu2.r_data_wire_3 ));
    InMux I__780 (
            .O(N__7062),
            .I(N__7059));
    LocalMux I__779 (
            .O(N__7059),
            .I(\uu2.un1_w_user_cr_5Z0Z_1 ));
    CascadeMux I__778 (
            .O(N__7056),
            .I(Lab_UT_L3_tx_data_2_0_cascade_));
    CascadeMux I__777 (
            .O(N__7053),
            .I(N__7049));
    InMux I__776 (
            .O(N__7052),
            .I(N__7044));
    InMux I__775 (
            .O(N__7049),
            .I(N__7044));
    LocalMux I__774 (
            .O(N__7044),
            .I(\uu2.un1_w_user_crZ0Z_5 ));
    InMux I__773 (
            .O(N__7041),
            .I(N__7038));
    LocalMux I__772 (
            .O(N__7038),
            .I(N__7034));
    InMux I__771 (
            .O(N__7037),
            .I(N__7031));
    Odrv4 I__770 (
            .O(N__7034),
            .I(Lab_UT_L3_tx_data_0_6));
    LocalMux I__769 (
            .O(N__7031),
            .I(Lab_UT_L3_tx_data_0_6));
    InMux I__768 (
            .O(N__7026),
            .I(N__7023));
    LocalMux I__767 (
            .O(N__7023),
            .I(\uu2.mem0.w_data_6 ));
    CascadeMux I__766 (
            .O(N__7020),
            .I(N__7016));
    InMux I__765 (
            .O(N__7019),
            .I(N__7011));
    InMux I__764 (
            .O(N__7016),
            .I(N__7008));
    InMux I__763 (
            .O(N__7015),
            .I(N__7003));
    InMux I__762 (
            .O(N__7014),
            .I(N__7003));
    LocalMux I__761 (
            .O(N__7011),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__760 (
            .O(N__7008),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__759 (
            .O(N__7003),
            .I(\uu2.w_addr_userZ0Z_8 ));
    CascadeMux I__758 (
            .O(N__6996),
            .I(N__6993));
    InMux I__757 (
            .O(N__6993),
            .I(N__6990));
    LocalMux I__756 (
            .O(N__6990),
            .I(\uu2.mem0.w_addr_8 ));
    InMux I__755 (
            .O(N__6987),
            .I(N__6984));
    LocalMux I__754 (
            .O(N__6984),
            .I(Lab_UT_L3_tx_data_2_0));
    CascadeMux I__753 (
            .O(N__6981),
            .I(N__6978));
    InMux I__752 (
            .O(N__6978),
            .I(N__6975));
    LocalMux I__751 (
            .O(N__6975),
            .I(\uu2.mem0.w_addr_1 ));
    InMux I__750 (
            .O(N__6972),
            .I(N__6969));
    LocalMux I__749 (
            .O(N__6969),
            .I(N__6963));
    InMux I__748 (
            .O(N__6968),
            .I(N__6958));
    InMux I__747 (
            .O(N__6967),
            .I(N__6958));
    InMux I__746 (
            .O(N__6966),
            .I(N__6955));
    Odrv4 I__745 (
            .O(N__6963),
            .I(L3_tx_data_2));
    LocalMux I__744 (
            .O(N__6958),
            .I(L3_tx_data_2));
    LocalMux I__743 (
            .O(N__6955),
            .I(L3_tx_data_2));
    InMux I__742 (
            .O(N__6948),
            .I(N__6945));
    LocalMux I__741 (
            .O(N__6945),
            .I(\uu2.mem0.w_data_2 ));
    InMux I__740 (
            .O(N__6942),
            .I(N__6936));
    InMux I__739 (
            .O(N__6941),
            .I(N__6936));
    LocalMux I__738 (
            .O(N__6936),
            .I(\uu2.un27_w_addr_user_0 ));
    InMux I__737 (
            .O(N__6933),
            .I(N__6928));
    InMux I__736 (
            .O(N__6932),
            .I(N__6925));
    InMux I__735 (
            .O(N__6931),
            .I(N__6922));
    LocalMux I__734 (
            .O(N__6928),
            .I(\Lab_UT.dspStr.cntZ0Z_0 ));
    LocalMux I__733 (
            .O(N__6925),
            .I(\Lab_UT.dspStr.cntZ0Z_0 ));
    LocalMux I__732 (
            .O(N__6922),
            .I(\Lab_UT.dspStr.cntZ0Z_0 ));
    InMux I__731 (
            .O(N__6915),
            .I(N__6912));
    LocalMux I__730 (
            .O(N__6912),
            .I(\uu2.un1_w_user_lfZ0Z_1 ));
    InMux I__729 (
            .O(N__6909),
            .I(N__6906));
    LocalMux I__728 (
            .O(N__6906),
            .I(\uu2.un1_w_user_lfZ0Z_3 ));
    InMux I__727 (
            .O(N__6903),
            .I(N__6900));
    LocalMux I__726 (
            .O(N__6900),
            .I(\uu2.un1_w_user_cr_0_0 ));
    InMux I__725 (
            .O(N__6897),
            .I(N__6894));
    LocalMux I__724 (
            .O(N__6894),
            .I(\uu2.un1_w_user_crZ0Z_2 ));
    InMux I__723 (
            .O(N__6891),
            .I(N__6888));
    LocalMux I__722 (
            .O(N__6888),
            .I(L3_tx_data_rdy));
    CascadeMux I__721 (
            .O(N__6885),
            .I(\uu2.un1_w_user_crZ0Z_2_cascade_ ));
    CascadeMux I__720 (
            .O(N__6882),
            .I(\uu2.un19_w_addr_userZ0Z_0_cascade_ ));
    InMux I__719 (
            .O(N__6879),
            .I(N__6873));
    InMux I__718 (
            .O(N__6878),
            .I(N__6873));
    LocalMux I__717 (
            .O(N__6873),
            .I(L3_tx_data_7));
    InMux I__716 (
            .O(N__6870),
            .I(N__6867));
    LocalMux I__715 (
            .O(N__6867),
            .I(N__6864));
    Span4Mux_h I__714 (
            .O(N__6864),
            .I(N__6861));
    Odrv4 I__713 (
            .O(N__6861),
            .I(\uu2.mem0.w_data_7 ));
    CascadeMux I__712 (
            .O(N__6858),
            .I(\Lab_UT.dspStr.cnt11_1_cascade_ ));
    InMux I__711 (
            .O(N__6855),
            .I(N__6851));
    CascadeMux I__710 (
            .O(N__6854),
            .I(N__6848));
    LocalMux I__709 (
            .O(N__6851),
            .I(N__6845));
    InMux I__708 (
            .O(N__6848),
            .I(N__6842));
    Odrv4 I__707 (
            .O(N__6845),
            .I(\Lab_UT.dspStr.cnt11_0_i ));
    LocalMux I__706 (
            .O(N__6842),
            .I(\Lab_UT.dspStr.cnt11_0_i ));
    IoInMux I__705 (
            .O(N__6837),
            .I(N__6834));
    LocalMux I__704 (
            .O(N__6834),
            .I(N__6831));
    IoSpan4Mux I__703 (
            .O(N__6831),
            .I(N__6828));
    Span4Mux_s2_h I__702 (
            .O(N__6828),
            .I(N__6825));
    Odrv4 I__701 (
            .O(N__6825),
            .I(\Lab_UT.secuu0.un11_l_count_i ));
    InMux I__700 (
            .O(N__6822),
            .I(N__6819));
    LocalMux I__699 (
            .O(N__6819),
            .I(Lab_UT_dspStr_un29_dOut_0));
    CascadeMux I__698 (
            .O(N__6816),
            .I(N__6811));
    CascadeMux I__697 (
            .O(N__6815),
            .I(N__6808));
    InMux I__696 (
            .O(N__6814),
            .I(N__6801));
    InMux I__695 (
            .O(N__6811),
            .I(N__6801));
    InMux I__694 (
            .O(N__6808),
            .I(N__6801));
    LocalMux I__693 (
            .O(N__6801),
            .I(\Lab_UT.secuu0.l_precountZ0Z_3 ));
    CascadeMux I__692 (
            .O(N__6798),
            .I(N__6793));
    InMux I__691 (
            .O(N__6797),
            .I(N__6785));
    InMux I__690 (
            .O(N__6796),
            .I(N__6785));
    InMux I__689 (
            .O(N__6793),
            .I(N__6785));
    InMux I__688 (
            .O(N__6792),
            .I(N__6782));
    LocalMux I__687 (
            .O(N__6785),
            .I(\Lab_UT.secuu0.l_countZ0Z_1 ));
    LocalMux I__686 (
            .O(N__6782),
            .I(\Lab_UT.secuu0.l_countZ0Z_1 ));
    InMux I__685 (
            .O(N__6777),
            .I(N__6762));
    InMux I__684 (
            .O(N__6776),
            .I(N__6762));
    InMux I__683 (
            .O(N__6775),
            .I(N__6762));
    InMux I__682 (
            .O(N__6774),
            .I(N__6762));
    InMux I__681 (
            .O(N__6773),
            .I(N__6762));
    LocalMux I__680 (
            .O(N__6762),
            .I(\Lab_UT.secuu0.l_precountZ0Z_1 ));
    InMux I__679 (
            .O(N__6759),
            .I(N__6753));
    InMux I__678 (
            .O(N__6758),
            .I(N__6748));
    InMux I__677 (
            .O(N__6757),
            .I(N__6748));
    InMux I__676 (
            .O(N__6756),
            .I(N__6745));
    LocalMux I__675 (
            .O(N__6753),
            .I(\Lab_UT.secuu0.l_countZ0Z_2 ));
    LocalMux I__674 (
            .O(N__6748),
            .I(\Lab_UT.secuu0.l_countZ0Z_2 ));
    LocalMux I__673 (
            .O(N__6745),
            .I(\Lab_UT.secuu0.l_countZ0Z_2 ));
    CascadeMux I__672 (
            .O(N__6738),
            .I(N__6732));
    InMux I__671 (
            .O(N__6737),
            .I(N__6723));
    InMux I__670 (
            .O(N__6736),
            .I(N__6723));
    InMux I__669 (
            .O(N__6735),
            .I(N__6723));
    InMux I__668 (
            .O(N__6732),
            .I(N__6723));
    LocalMux I__667 (
            .O(N__6723),
            .I(\Lab_UT.secuu0.l_precountZ0Z_2 ));
    InMux I__666 (
            .O(N__6720),
            .I(N__6707));
    InMux I__665 (
            .O(N__6719),
            .I(N__6707));
    InMux I__664 (
            .O(N__6718),
            .I(N__6707));
    InMux I__663 (
            .O(N__6717),
            .I(N__6707));
    InMux I__662 (
            .O(N__6716),
            .I(N__6704));
    LocalMux I__661 (
            .O(N__6707),
            .I(\Lab_UT.secuu0.l_countZ0Z_0 ));
    LocalMux I__660 (
            .O(N__6704),
            .I(\Lab_UT.secuu0.l_countZ0Z_0 ));
    CascadeMux I__659 (
            .O(N__6699),
            .I(\Lab_UT.secuu0.un4_l_count_14_cascade_ ));
    InMux I__658 (
            .O(N__6696),
            .I(N__6691));
    InMux I__657 (
            .O(N__6695),
            .I(N__6686));
    InMux I__656 (
            .O(N__6694),
            .I(N__6686));
    LocalMux I__655 (
            .O(N__6691),
            .I(N__6680));
    LocalMux I__654 (
            .O(N__6686),
            .I(N__6680));
    InMux I__653 (
            .O(N__6685),
            .I(N__6677));
    Odrv4 I__652 (
            .O(N__6680),
            .I(\Lab_UT.secuu0.un4_l_count_0_8 ));
    LocalMux I__651 (
            .O(N__6677),
            .I(\Lab_UT.secuu0.un4_l_count_0_8 ));
    InMux I__650 (
            .O(N__6672),
            .I(N__6669));
    LocalMux I__649 (
            .O(N__6669),
            .I(\Lab_UT.secuu0.un4_l_count_12 ));
    InMux I__648 (
            .O(N__6666),
            .I(N__6663));
    LocalMux I__647 (
            .O(N__6663),
            .I(\Lab_UT.secuu0.un4_l_count_13 ));
    CascadeMux I__646 (
            .O(N__6660),
            .I(\Lab_UT.secuu0.un4_l_count_18_cascade_ ));
    CascadeMux I__645 (
            .O(N__6657),
            .I(N__6654));
    InMux I__644 (
            .O(N__6654),
            .I(N__6651));
    LocalMux I__643 (
            .O(N__6651),
            .I(N__6648));
    Odrv4 I__642 (
            .O(N__6648),
            .I(\Lab_UT.secuu0.un230_ci_1 ));
    CascadeMux I__641 (
            .O(N__6645),
            .I(N__6639));
    InMux I__640 (
            .O(N__6644),
            .I(N__6636));
    InMux I__639 (
            .O(N__6643),
            .I(N__6633));
    InMux I__638 (
            .O(N__6642),
            .I(N__6627));
    InMux I__637 (
            .O(N__6639),
            .I(N__6627));
    LocalMux I__636 (
            .O(N__6636),
            .I(N__6624));
    LocalMux I__635 (
            .O(N__6633),
            .I(N__6621));
    InMux I__634 (
            .O(N__6632),
            .I(N__6618));
    LocalMux I__633 (
            .O(N__6627),
            .I(\Lab_UT.secuu0.un109_ci ));
    Odrv4 I__632 (
            .O(N__6624),
            .I(\Lab_UT.secuu0.un109_ci ));
    Odrv4 I__631 (
            .O(N__6621),
            .I(\Lab_UT.secuu0.un109_ci ));
    LocalMux I__630 (
            .O(N__6618),
            .I(\Lab_UT.secuu0.un109_ci ));
    CascadeMux I__629 (
            .O(N__6609),
            .I(\Lab_UT.secuu0.un197_ci_9_cascade_ ));
    InMux I__628 (
            .O(N__6606),
            .I(N__6600));
    InMux I__627 (
            .O(N__6605),
            .I(N__6593));
    InMux I__626 (
            .O(N__6604),
            .I(N__6593));
    InMux I__625 (
            .O(N__6603),
            .I(N__6593));
    LocalMux I__624 (
            .O(N__6600),
            .I(\Lab_UT.secuu0.l_countZ0Z_14 ));
    LocalMux I__623 (
            .O(N__6593),
            .I(\Lab_UT.secuu0.l_countZ0Z_14 ));
    CascadeMux I__622 (
            .O(N__6588),
            .I(N__6583));
    CascadeMux I__621 (
            .O(N__6587),
            .I(N__6580));
    InMux I__620 (
            .O(N__6586),
            .I(N__6573));
    InMux I__619 (
            .O(N__6583),
            .I(N__6573));
    InMux I__618 (
            .O(N__6580),
            .I(N__6573));
    LocalMux I__617 (
            .O(N__6573),
            .I(\Lab_UT.secuu0.l_countZ0Z_15 ));
    CascadeMux I__616 (
            .O(N__6570),
            .I(N__6565));
    InMux I__615 (
            .O(N__6569),
            .I(N__6561));
    InMux I__614 (
            .O(N__6568),
            .I(N__6558));
    InMux I__613 (
            .O(N__6565),
            .I(N__6553));
    InMux I__612 (
            .O(N__6564),
            .I(N__6553));
    LocalMux I__611 (
            .O(N__6561),
            .I(\Lab_UT.secuu0.l_countZ0Z_4 ));
    LocalMux I__610 (
            .O(N__6558),
            .I(\Lab_UT.secuu0.l_countZ0Z_4 ));
    LocalMux I__609 (
            .O(N__6553),
            .I(\Lab_UT.secuu0.l_countZ0Z_4 ));
    InMux I__608 (
            .O(N__6546),
            .I(N__6541));
    InMux I__607 (
            .O(N__6545),
            .I(N__6538));
    InMux I__606 (
            .O(N__6544),
            .I(N__6535));
    LocalMux I__605 (
            .O(N__6541),
            .I(N__6532));
    LocalMux I__604 (
            .O(N__6538),
            .I(\Lab_UT.secuu0.l_countZ0Z_5 ));
    LocalMux I__603 (
            .O(N__6535),
            .I(\Lab_UT.secuu0.l_countZ0Z_5 ));
    Odrv4 I__602 (
            .O(N__6532),
            .I(\Lab_UT.secuu0.l_countZ0Z_5 ));
    InMux I__601 (
            .O(N__6525),
            .I(N__6522));
    LocalMux I__600 (
            .O(N__6522),
            .I(uart_RXD));
    CascadeMux I__599 (
            .O(N__6519),
            .I(\uu2.un447_ci_3_cascade_ ));
    InMux I__598 (
            .O(N__6516),
            .I(N__6513));
    LocalMux I__597 (
            .O(N__6513),
            .I(\uu2.o_adder_vbuf_w_addr_user_7 ));
    CascadeMux I__596 (
            .O(N__6510),
            .I(N__6507));
    InMux I__595 (
            .O(N__6507),
            .I(N__6504));
    LocalMux I__594 (
            .O(N__6504),
            .I(N__6501));
    Span4Mux_v I__593 (
            .O(N__6501),
            .I(N__6498));
    Odrv4 I__592 (
            .O(N__6498),
            .I(\uu2.mem0.w_addr_6 ));
    CascadeMux I__591 (
            .O(N__6495),
            .I(N__6492));
    InMux I__590 (
            .O(N__6492),
            .I(N__6489));
    LocalMux I__589 (
            .O(N__6489),
            .I(N__6486));
    Span4Mux_h I__588 (
            .O(N__6486),
            .I(N__6483));
    Odrv4 I__587 (
            .O(N__6483),
            .I(\uu2.mem0.w_addr_7 ));
    InMux I__586 (
            .O(N__6480),
            .I(N__6473));
    InMux I__585 (
            .O(N__6479),
            .I(N__6464));
    InMux I__584 (
            .O(N__6478),
            .I(N__6464));
    InMux I__583 (
            .O(N__6477),
            .I(N__6464));
    InMux I__582 (
            .O(N__6476),
            .I(N__6464));
    LocalMux I__581 (
            .O(N__6473),
            .I(\uu2.w_addr_userZ0Z_6 ));
    LocalMux I__580 (
            .O(N__6464),
            .I(\uu2.w_addr_userZ0Z_6 ));
    InMux I__579 (
            .O(N__6459),
            .I(N__6452));
    InMux I__578 (
            .O(N__6458),
            .I(N__6447));
    InMux I__577 (
            .O(N__6457),
            .I(N__6447));
    InMux I__576 (
            .O(N__6456),
            .I(N__6442));
    InMux I__575 (
            .O(N__6455),
            .I(N__6442));
    LocalMux I__574 (
            .O(N__6452),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__573 (
            .O(N__6447),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__572 (
            .O(N__6442),
            .I(\uu2.w_addr_userZ0Z_7 ));
    CascadeMux I__571 (
            .O(N__6435),
            .I(N__6432));
    InMux I__570 (
            .O(N__6432),
            .I(N__6428));
    InMux I__569 (
            .O(N__6431),
            .I(N__6425));
    LocalMux I__568 (
            .O(N__6428),
            .I(\uu2.un447_ci_3 ));
    LocalMux I__567 (
            .O(N__6425),
            .I(\uu2.un447_ci_3 ));
    CascadeMux I__566 (
            .O(N__6420),
            .I(\uu2.vbuf_w_addr_user.un469_ci_0_cascade_ ));
    CascadeMux I__565 (
            .O(N__6417),
            .I(N__6414));
    InMux I__564 (
            .O(N__6414),
            .I(N__6411));
    LocalMux I__563 (
            .O(N__6411),
            .I(\uu2.o_adder_vbuf_w_addr_user_8 ));
    InMux I__562 (
            .O(N__6408),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_2 ));
    InMux I__561 (
            .O(N__6405),
            .I(N__6402));
    LocalMux I__560 (
            .O(N__6402),
            .I(N__6399));
    Odrv4 I__559 (
            .O(N__6399),
            .I(\uu2.un1_w_user_lfZ0Z_4 ));
    CascadeMux I__558 (
            .O(N__6396),
            .I(L3_tx_data_0_cascade_));
    InMux I__557 (
            .O(N__6393),
            .I(N__6390));
    LocalMux I__556 (
            .O(N__6390),
            .I(\uu2.un1_w_user_lf_0 ));
    CascadeMux I__555 (
            .O(N__6387),
            .I(\uu2.un1_w_user_lf_0_cascade_ ));
    CascadeMux I__554 (
            .O(N__6384),
            .I(Lab_UT_L3_tx_data_0_4_cascade_));
    CascadeMux I__553 (
            .O(N__6381),
            .I(Lab_UT_dspStr_un29_dOut_0_cascade_));
    InMux I__552 (
            .O(N__6378),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_0 ));
    InMux I__551 (
            .O(N__6375),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_1 ));
    CascadeMux I__550 (
            .O(N__6372),
            .I(N__6369));
    InMux I__549 (
            .O(N__6369),
            .I(N__6366));
    LocalMux I__548 (
            .O(N__6366),
            .I(\Lab_UT.secuu0.un142_ci_0 ));
    CascadeMux I__547 (
            .O(N__6363),
            .I(N__6359));
    InMux I__546 (
            .O(N__6362),
            .I(N__6354));
    InMux I__545 (
            .O(N__6359),
            .I(N__6354));
    LocalMux I__544 (
            .O(N__6354),
            .I(\Lab_UT.secuu0.un131_ci_3 ));
    InMux I__543 (
            .O(N__6351),
            .I(N__6348));
    LocalMux I__542 (
            .O(N__6348),
            .I(\Lab_UT.secuu0.un87_ci ));
    CascadeMux I__541 (
            .O(N__6345),
            .I(\Lab_UT.secuu0.un87_ci_cascade_ ));
    CascadeMux I__540 (
            .O(N__6342),
            .I(\Lab_UT.secuu0.un131_ci_3_cascade_ ));
    IoInMux I__539 (
            .O(N__6339),
            .I(N__6336));
    LocalMux I__538 (
            .O(N__6336),
            .I(N__6333));
    IoSpan4Mux I__537 (
            .O(N__6333),
            .I(N__6330));
    Odrv4 I__536 (
            .O(N__6330),
            .I(clk_in_c));
    INV \INVuu2.w_addr_displaying_0C  (
            .O(\INVuu2.w_addr_displaying_0C_net ),
            .I(N__13494));
    INV \INVuu2.w_addr_displaying_2_rep1C  (
            .O(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .I(N__13499));
    INV \INVuu2.w_addr_displaying_0_rep1C  (
            .O(\INVuu2.w_addr_displaying_0_rep1C_net ),
            .I(N__13504));
    INV \INVuu2.w_addr_displaying_4_rep1C  (
            .O(\INVuu2.w_addr_displaying_4_rep1C_net ),
            .I(N__13520));
    INV \INVuu2.w_addr_displaying_fast_3C  (
            .O(\INVuu2.w_addr_displaying_fast_3C_net ),
            .I(N__13498));
    INV \INVuu2.w_addr_displaying_6_rep1C  (
            .O(\INVuu2.w_addr_displaying_6_rep1C_net ),
            .I(N__13503));
    INV \INVuu2.w_addr_displaying_6C  (
            .O(\INVuu2.w_addr_displaying_6C_net ),
            .I(N__13512));
    INV \INVuu2.w_addr_displaying_2C  (
            .O(\INVuu2.w_addr_displaying_2C_net ),
            .I(N__13484));
    INV \INVuu2.w_addr_displaying_4C  (
            .O(\INVuu2.w_addr_displaying_4C_net ),
            .I(N__13492));
    INV \INVuu2.w_addr_displaying_fast_4C  (
            .O(\INVuu2.w_addr_displaying_fast_4C_net ),
            .I(N__13497));
    INV \INVuu2.w_addr_displaying_5C  (
            .O(\INVuu2.w_addr_displaying_5C_net ),
            .I(N__13483));
    INV \INVuu2.w_addr_displaying_1C  (
            .O(\INVuu2.w_addr_displaying_1C_net ),
            .I(N__13491));
    INV \INVuu2.w_addr_user_3C  (
            .O(\INVuu2.w_addr_user_3C_net ),
            .I(N__13507));
    INV \INVuu2.w_addr_user_4C  (
            .O(\INVuu2.w_addr_user_4C_net ),
            .I(N__13515));
    defparam IN_MUX_bfv_7_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_2_0_));
    defparam IN_MUX_bfv_6_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_1_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_8_0_));
    ICE_GB \latticehx1k_pll_inst.PLLOUTCORE_derived_clock_RNIALC1  (
            .USERSIGNALTOGLOBALBUFFER(N__8142),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB \Lab_UT.secuu0.delay_line_RNILBAI7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__6837),
            .GLOBALBUFFEROUTPUT(\Lab_UT.secuu0.un11_l_count_i_g ));
    GND GND (
            .Y(GNDG0));
    ICE_GB \resetGen.rst_RNI4PQ1  (
            .USERSIGNALTOGLOBALBUFFER(N__10931),
            .GLOBALBUFFEROUTPUT(rst_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_5_LC_1_3_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_5_LC_1_3_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_5_LC_1_3_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \Lab_UT.secuu0.l_count_5_LC_1_3_0  (
            .in0(N__6643),
            .in1(N__6545),
            .in2(_gnd_net_),
            .in3(N__6569),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13548),
            .ce(N__7583),
            .sr(N__15898));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_3_LC_1_4_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_3_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_3_LC_1_4_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_3_LC_1_4_1  (
            .in0(_gnd_net_),
            .in1(N__6544),
            .in2(_gnd_net_),
            .in3(N__6568),
            .lcout(\Lab_UT.secuu0.un131_ci_3 ),
            .ltout(\Lab_UT.secuu0.un131_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_7__un142_ci_0_LC_1_4_2 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_7__un142_ci_0_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_7__un142_ci_0_LC_1_4_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_7__un142_ci_0_LC_1_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6342),
            .in3(N__7343),
            .lcout(\Lab_UT.secuu0.un142_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_15__un230_ci_1_LC_1_4_7 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_15__un230_ci_1_LC_1_4_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_15__un230_ci_1_LC_1_4_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_15__un230_ci_1_LC_1_4_7  (
            .in0(N__6696),
            .in1(N__7726),
            .in2(_gnd_net_),
            .in3(N__6606),
            .lcout(\Lab_UT.secuu0.un230_ci_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_3_LC_1_5_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_3_LC_1_5_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_3_LC_1_5_3 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \Lab_UT.secuu0.l_count_3_LC_1_5_3  (
            .in0(N__6351),
            .in1(N__6759),
            .in2(N__7395),
            .in3(N__11044),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13545),
            .ce(N__7582),
            .sr(N__15896));
    defparam \Lab_UT.secuu0.l_count_7_LC_1_5_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_7_LC_1_5_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_7_LC_1_5_4 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Lab_UT.secuu0.l_count_7_LC_1_5_4  (
            .in0(N__11043),
            .in1(N__6642),
            .in2(N__6372),
            .in3(N__7412),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13545),
            .ce(N__7582),
            .sr(N__15896));
    defparam \Lab_UT.secuu0.l_count_6_LC_1_5_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_6_LC_1_5_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_6_LC_1_5_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \Lab_UT.secuu0.l_count_6_LC_1_5_5  (
            .in0(N__7342),
            .in1(N__6362),
            .in2(N__6645),
            .in3(N__11042),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13545),
            .ce(N__7582),
            .sr(N__15896));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_8_LC_1_5_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_8_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_8_LC_1_5_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_8_LC_1_5_6  (
            .in0(N__6632),
            .in1(N__7341),
            .in2(N__6363),
            .in3(N__7411),
            .lcout(\Lab_UT.secuu0.un153_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_6_LC_1_6_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_6_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_6_LC_1_6_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_6_LC_1_6_0  (
            .in0(N__6757),
            .in1(N__6717),
            .in2(N__6798),
            .in3(N__7390),
            .lcout(\Lab_UT.secuu0.un109_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_1_LC_1_6_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_1_LC_1_6_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_1_LC_1_6_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.secuu0.l_count_1_LC_1_6_1  (
            .in0(N__6720),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6797),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13541),
            .ce(N__7581),
            .sr(N__15895));
    defparam \Lab_UT.secuu0.l_count_0_LC_1_6_2 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_0_LC_1_6_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_0_LC_1_6_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.secuu0.l_count_0_LC_1_6_2  (
            .in0(_gnd_net_),
            .in1(N__6719),
            .in2(_gnd_net_),
            .in3(N__11045),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13541),
            .ce(N__7581),
            .sr(N__15895));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_1_LC_1_6_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_1_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_1_LC_1_6_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_1_LC_1_6_3  (
            .in0(N__6718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6796),
            .lcout(\Lab_UT.secuu0.un87_ci ),
            .ltout(\Lab_UT.secuu0.un87_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_2_LC_1_6_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_2_LC_1_6_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_2_LC_1_6_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \Lab_UT.secuu0.l_count_2_LC_1_6_4  (
            .in0(N__6758),
            .in1(_gnd_net_),
            .in2(N__6345),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13541),
            .ce(N__7581),
            .sr(N__15895));
    defparam \Lab_UT.secuu0.l_count_RNIFM2M_13_LC_1_6_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNIFM2M_13_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNIFM2M_13_LC_1_6_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNIFM2M_13_LC_1_6_6  (
            .in0(N__7604),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7704),
            .lcout(\Lab_UT.secuu0.un4_l_count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNIMHJI1_2_LC_1_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNIMHJI1_2_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNIMHJI1_2_LC_1_7_0 .LUT_INIT=16'b1010011111100111;
    LogicCell40 \Lab_UT.dspStr.cnt_RNIMHJI1_2_LC_1_7_0  (
            .in0(N__8562),
            .in1(N__8728),
            .in2(N__8666),
            .in3(N__8842),
            .lcout(),
            .ltout(Lab_UT_L3_tx_data_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_4_LC_1_7_1 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_4_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_4_LC_1_7_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \uu2.un1_w_user_lf_4_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6384),
            .in3(N__6966),
            .lcout(\uu2.un1_w_user_lfZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNIKFJI1_2_LC_1_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNIKFJI1_2_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNIKFJI1_2_LC_1_7_2 .LUT_INIT=16'b1110000110100001;
    LogicCell40 \Lab_UT.dspStr.cnt_RNIKFJI1_2_LC_1_7_2  (
            .in0(N__8561),
            .in1(N__8726),
            .in2(N__8665),
            .in3(N__10297),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.Lab3U00.q_esr_2_LC_1_7_4 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_2_LC_1_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_2_LC_1_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_2_LC_1_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9666),
            .lcout(\Lab_UT.rx_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13533),
            .ce(N__9090),
            .sr(N__15873));
    defparam \Lab_UT.dspStr.cnt_RNI57RQ_2_LC_1_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNI57RQ_2_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNI57RQ_2_LC_1_7_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dspStr.cnt_RNI57RQ_2_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(N__8642),
            .in2(_gnd_net_),
            .in3(N__8560),
            .lcout(Lab_UT_dspStr_un29_dOut_0),
            .ltout(Lab_UT_dspStr_un29_dOut_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_0_LC_1_7_6 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_0_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_0_LC_1_7_6 .LUT_INIT=16'b0011111101111111;
    LogicCell40 \uu2.un1_w_user_cr_0_LC_1_7_6  (
            .in0(N__8841),
            .in1(N__8727),
            .in2(N__6381),
            .in3(N__8774),
            .lcout(\uu2.un1_w_user_cr_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_0_LC_1_8_0 .C_ON=1'b1;
    defparam \Lab_UT.dspStr.cnt_0_LC_1_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_0_LC_1_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.dspStr.cnt_0_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__6932),
            .in2(N__6854),
            .in3(N__6855),
            .lcout(\Lab_UT.dspStr.cntZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(\Lab_UT.dspStr.un1_cnt_3_cry_0 ),
            .clk(N__13528),
            .ce(),
            .sr(N__15872));
    defparam \Lab_UT.dspStr.cnt_1_LC_1_8_1 .C_ON=1'b1;
    defparam \Lab_UT.dspStr.cnt_1_LC_1_8_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_1_LC_1_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.dspStr.cnt_1_LC_1_8_1  (
            .in0(_gnd_net_),
            .in1(N__8742),
            .in2(_gnd_net_),
            .in3(N__6378),
            .lcout(Lab_UT_dspStr_cnt_1),
            .ltout(),
            .carryin(\Lab_UT.dspStr.un1_cnt_3_cry_0 ),
            .carryout(\Lab_UT.dspStr.un1_cnt_3_cry_1 ),
            .clk(N__13528),
            .ce(),
            .sr(N__15872));
    defparam \Lab_UT.dspStr.cnt_2_LC_1_8_2 .C_ON=1'b1;
    defparam \Lab_UT.dspStr.cnt_2_LC_1_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_2_LC_1_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.dspStr.cnt_2_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(N__8574),
            .in2(_gnd_net_),
            .in3(N__6375),
            .lcout(Lab_UT_dspStr_cnt_2),
            .ltout(),
            .carryin(\Lab_UT.dspStr.un1_cnt_3_cry_1 ),
            .carryout(\Lab_UT.dspStr.un1_cnt_3_cry_2 ),
            .clk(N__13528),
            .ce(),
            .sr(N__15872));
    defparam \Lab_UT.dspStr.cnt_3_LC_1_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_3_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_3_LC_1_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.dspStr.cnt_3_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(N__8664),
            .in2(_gnd_net_),
            .in3(N__6408),
            .lcout(Lab_UT_dspStr_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13528),
            .ce(),
            .sr(N__15872));
    defparam \uu2.w_addr_user_RNIKHHEL_2_LC_1_9_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIKHHEL_2_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIKHHEL_2_LC_1_9_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \uu2.w_addr_user_RNIKHHEL_2_LC_1_9_0  (
            .in0(N__10938),
            .in1(N__6942),
            .in2(_gnd_net_),
            .in3(N__6393),
            .lcout(\uu2.w_addr_user_RNIKHHELZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNIIDJI1_0_2_LC_1_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNIIDJI1_0_2_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNIIDJI1_0_2_LC_1_9_4 .LUT_INIT=16'b1110111010100010;
    LogicCell40 \Lab_UT.dspStr.cnt_RNIIDJI1_0_2_LC_1_9_4  (
            .in0(N__8741),
            .in1(N__8660),
            .in2(N__10370),
            .in3(N__8570),
            .lcout(),
            .ltout(L3_tx_data_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_LC_1_9_5 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_LC_1_9_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uu2.un1_w_user_lf_LC_1_9_5  (
            .in0(N__8162),
            .in1(N__6405),
            .in2(N__6396),
            .in3(N__6909),
            .lcout(\uu2.un1_w_user_lf_0 ),
            .ltout(\uu2.un1_w_user_lf_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNILJEE01_2_LC_1_9_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNILJEE01_2_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNILJEE01_2_LC_1_9_6 .LUT_INIT=16'b1111111111110011;
    LogicCell40 \uu2.w_addr_user_RNILJEE01_2_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(N__6941),
            .in2(N__6387),
            .in3(N__12399),
            .lcout(\uu2.un27_w_addr_user_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_4_LC_1_10_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_4_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_4_LC_1_10_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.w_addr_user_4_LC_1_10_0  (
            .in0(N__7099),
            .in1(N__9371),
            .in2(_gnd_net_),
            .in3(N__7194),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_4C_net ),
            .ce(),
            .sr(N__7160));
    defparam \uu2.w_addr_user_8_LC_1_10_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_8_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_8_LC_1_10_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \uu2.w_addr_user_8_LC_1_10_1  (
            .in0(N__7196),
            .in1(_gnd_net_),
            .in2(N__6417),
            .in3(N__7019),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_4C_net ),
            .ce(),
            .sr(N__7160));
    defparam \uu2.w_addr_user_7_LC_1_10_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_7_LC_1_10_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_7_LC_1_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.w_addr_user_7_LC_1_10_4  (
            .in0(N__6516),
            .in1(N__6459),
            .in2(_gnd_net_),
            .in3(N__7195),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_4C_net ),
            .ce(),
            .sr(N__7160));
    defparam \uu2.w_addr_user_6_LC_1_10_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_6_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_6_LC_1_10_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_6_LC_1_10_7  (
            .in0(N__7197),
            .in1(N__7100),
            .in2(N__6435),
            .in3(N__6480),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_4C_net ),
            .ce(),
            .sr(N__7160));
    defparam \buart.Z_rx.hh_0_LC_1_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_1_11_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.hh_0_LC_1_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6525),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13506),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un447_ci_3_LC_1_11_1 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un447_ci_3_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un447_ci_3_LC_1_11_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_6__un447_ci_3_LC_1_11_1  (
            .in0(N__9322),
            .in1(N__9370),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.un447_ci_3 ),
            .ltout(\uu2.un447_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.result_1_7_LC_1_11_2 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.result_1_7_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.result_1_7_LC_1_11_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.vbuf_w_addr_user.result_1_7_LC_1_11_2  (
            .in0(N__6479),
            .in1(N__7094),
            .in2(N__6519),
            .in3(N__6458),
            .lcout(\uu2.o_adder_vbuf_w_addr_user_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_1_11_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_1_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_1_11_3  (
            .in0(N__12460),
            .in1(N__6477),
            .in2(_gnd_net_),
            .in3(N__12231),
            .lcout(\uu2.mem0.w_addr_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_1_11_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_1_11_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_1_11_4  (
            .in0(N__6456),
            .in1(N__12461),
            .in2(_gnd_net_),
            .in3(N__16290),
            .lcout(\uu2.mem0.w_addr_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIOGH7_8_LC_1_11_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIOGH7_8_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIOGH7_8_LC_1_11_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uu2.w_addr_user_RNIOGH7_8_LC_1_11_5  (
            .in0(N__7014),
            .in1(N__6455),
            .in2(_gnd_net_),
            .in3(N__6476),
            .lcout(\uu2.un2_w_addr_user_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un469_ci_0_LC_1_11_6 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un469_ci_0_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un469_ci_0_LC_1_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_8__un469_ci_0_LC_1_11_6  (
            .in0(N__6478),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6457),
            .lcout(),
            .ltout(\uu2.vbuf_w_addr_user.un469_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.result_1_8_LC_1_11_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.result_1_8_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.result_1_8_LC_1_11_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.vbuf_w_addr_user.result_1_8_LC_1_11_7  (
            .in0(N__7015),
            .in1(N__6431),
            .in2(N__6420),
            .in3(N__7095),
            .lcout(\uu2.o_adder_vbuf_w_addr_user_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_9_LC_2_3_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_9_LC_2_3_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_9_LC_2_3_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \Lab_UT.secuu0.l_count_9_LC_2_3_0  (
            .in0(N__7671),
            .in1(N__7494),
            .in2(_gnd_net_),
            .in3(N__7444),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13547),
            .ce(N__7586),
            .sr(N__15901));
    defparam \Lab_UT.secuu0.l_count_10_LC_2_4_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_10_LC_2_4_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_10_LC_2_4_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \Lab_UT.secuu0.l_count_10_LC_2_4_0  (
            .in0(N__7440),
            .in1(N__7517),
            .in2(N__7670),
            .in3(N__7489),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13546),
            .ce(N__7584),
            .sr(N__15899));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_16__un241_ci_2_LC_2_4_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_16__un241_ci_2_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_16__un241_ci_2_LC_2_4_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_16__un241_ci_2_LC_2_4_1  (
            .in0(N__6604),
            .in1(N__7720),
            .in2(N__6588),
            .in3(N__6694),
            .lcout(\Lab_UT.secuu0.un241_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_15_LC_2_4_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_15_LC_2_4_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_15_LC_2_4_3 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \Lab_UT.secuu0.l_count_15_LC_2_4_3  (
            .in0(N__6586),
            .in1(N__7646),
            .in2(N__6657),
            .in3(N__11040),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13546),
            .ce(N__7584),
            .sr(N__15899));
    defparam \Lab_UT.secuu0.l_count_4_LC_2_4_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_4_LC_2_4_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_4_LC_2_4_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \Lab_UT.secuu0.l_count_4_LC_2_4_4  (
            .in0(N__11041),
            .in1(_gnd_net_),
            .in2(N__6570),
            .in3(N__6644),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13546),
            .ce(N__7584),
            .sr(N__15899));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_12__un197_ci_9_LC_2_4_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_12__un197_ci_9_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_12__un197_ci_9_LC_2_4_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_12__un197_ci_9_LC_2_4_5  (
            .in0(N__7516),
            .in1(N__7439),
            .in2(N__7371),
            .in3(N__7488),
            .lcout(\Lab_UT.secuu0.un197_ci_9 ),
            .ltout(\Lab_UT.secuu0.un197_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_14_LC_2_4_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_14_LC_2_4_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_14_LC_2_4_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \Lab_UT.secuu0.l_count_14_LC_2_4_6  (
            .in0(N__6695),
            .in1(N__7674),
            .in2(N__6609),
            .in3(N__6605),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13546),
            .ce(N__7584),
            .sr(N__15899));
    defparam \Lab_UT.secuu0.l_count_RNIGLN81_15_LC_2_4_7 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNIGLN81_15_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNIGLN81_15_LC_2_4_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNIGLN81_15_LC_2_4_7  (
            .in0(N__6603),
            .in1(N__7515),
            .in2(N__6587),
            .in3(N__6564),
            .lcout(\Lab_UT.secuu0.un4_l_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.delay_line_0_LC_2_5_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.delay_line_0_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.delay_line_0_LC_2_5_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.delay_line_0_LC_2_5_0  (
            .in0(N__6774),
            .in1(N__7555),
            .in2(N__6816),
            .in3(N__6735),
            .lcout(\Lab_UT.secuu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13542),
            .ce(),
            .sr(N__15897));
    defparam \Lab_UT.secuu0.l_precount_3_LC_2_5_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_precount_3_LC_2_5_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_precount_3_LC_2_5_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \Lab_UT.secuu0.l_precount_3_LC_2_5_1  (
            .in0(N__6737),
            .in1(N__6814),
            .in2(N__7560),
            .in3(N__6777),
            .lcout(\Lab_UT.secuu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13542),
            .ce(),
            .sr(N__15897));
    defparam \Lab_UT.secuu0.l_count_RNI8TM21_5_LC_2_5_2 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNI8TM21_5_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNI8TM21_5_LC_2_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.secuu0.l_count_RNI8TM21_5_LC_2_5_2  (
            .in0(N__6773),
            .in1(N__6546),
            .in2(N__6815),
            .in3(N__6792),
            .lcout(\Lab_UT.secuu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_precount_1_LC_2_5_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_precount_1_LC_2_5_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_precount_1_LC_2_5_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.secuu0.l_precount_1_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(N__7554),
            .in2(_gnd_net_),
            .in3(N__6775),
            .lcout(\Lab_UT.secuu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13542),
            .ce(),
            .sr(N__15897));
    defparam \Lab_UT.secuu0.l_precount_2_LC_2_5_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_precount_2_LC_2_5_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_precount_2_LC_2_5_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \Lab_UT.secuu0.l_precount_2_LC_2_5_4  (
            .in0(N__6776),
            .in1(N__7556),
            .in2(_gnd_net_),
            .in3(N__6736),
            .lcout(\Lab_UT.secuu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13542),
            .ce(),
            .sr(N__15897));
    defparam \Lab_UT.secuu0.l_count_RNI3II01_2_LC_2_5_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNI3II01_2_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNI3II01_2_LC_2_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.secuu0.l_count_RNI3II01_2_LC_2_5_5  (
            .in0(N__7493),
            .in1(N__6756),
            .in2(N__6738),
            .in3(N__6716),
            .lcout(),
            .ltout(\Lab_UT.secuu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_RNIOIEB2_16_LC_2_5_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNIOIEB2_16_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNIOIEB2_16_LC_2_5_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNIOIEB2_16_LC_2_5_6  (
            .in0(N__7553),
            .in1(N__7263),
            .in2(N__6699),
            .in3(N__6685),
            .lcout(),
            .ltout(\Lab_UT.secuu0.un4_l_count_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_RNI82GM6_5_LC_2_5_7 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNI82GM6_5_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNI82GM6_5_LC_2_5_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNI82GM6_5_LC_2_5_7  (
            .in0(N__6672),
            .in1(N__6666),
            .in2(N__6660),
            .in3(N__7320),
            .lcout(\Lab_UT.secuu0.un4_l_count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.Lab3U00.q_esr_0_LC_2_6_0 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_0_LC_2_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_0_LC_2_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_0_LC_2_6_0  (
            .in0(N__13599),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.rx_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13534),
            .ce(N__9083),
            .sr(N__15875));
    defparam \Lab_UT.Lab3U00.q_esr_3_LC_2_6_1 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_3_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_3_LC_2_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_3_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9618),
            .lcout(Lab_UT_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13534),
            .ce(N__9083),
            .sr(N__15875));
    defparam \Lab_UT.Lab3U00.q_esr_5_LC_2_6_2 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_5_LC_2_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_5_LC_2_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_5_LC_2_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8499),
            .lcout(Lab_UT_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13534),
            .ce(N__9083),
            .sr(N__15875));
    defparam \Lab_UT.Lab3U00.q_esr_6_LC_2_6_3 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_6_LC_2_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_6_LC_2_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_6_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9690),
            .lcout(Lab_UT_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13534),
            .ce(N__9083),
            .sr(N__15875));
    defparam \Lab_UT.Lab3U00.q_esr_7_LC_2_6_4 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_7_LC_2_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_7_LC_2_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_7_LC_2_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9717),
            .lcout(Lab_UT_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13534),
            .ce(N__9083),
            .sr(N__15875));
    defparam \Lab_UT.Lab3U00.q_esr_4_LC_2_6_5 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_4_LC_2_6_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_4_LC_2_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_4_LC_2_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9642),
            .lcout(Lab_UT_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13534),
            .ce(N__9083),
            .sr(N__15875));
    defparam \Lab_UT.dspStr.cnt_RNI11B71_2_LC_2_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNI11B71_2_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNI11B71_2_LC_2_7_1 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \Lab_UT.dspStr.cnt_RNI11B71_2_LC_2_7_1  (
            .in0(N__16546),
            .in1(N__8654),
            .in2(N__13344),
            .in3(N__8565),
            .lcout(),
            .ltout(\Lab_UT.dspStr.cnt11_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNI24622_0_LC_2_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNI24622_0_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNI24622_0_LC_2_7_2 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \Lab_UT.dspStr.cnt_RNI24622_0_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__6931),
            .in2(N__6858),
            .in3(N__8724),
            .lcout(\Lab_UT.dspStr.cnt11_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.delay_line_RNILBAI7_1_LC_2_7_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.delay_line_RNILBAI7_1_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.delay_line_RNILBAI7_1_LC_2_7_3 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \Lab_UT.secuu0.delay_line_RNILBAI7_1_LC_2_7_3  (
            .in0(N__10974),
            .in1(N__10988),
            .in2(_gnd_net_),
            .in3(N__11052),
            .lcout(\Lab_UT.secuu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_1_LC_2_7_4 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_1_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_1_LC_2_7_4 .LUT_INIT=16'b0011011111111111;
    LogicCell40 \uu2.un1_w_user_lf_1_LC_2_7_4  (
            .in0(N__8772),
            .in1(N__8723),
            .in2(N__10225),
            .in3(N__6822),
            .lcout(\uu2.un1_w_user_lfZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_2_7_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_2_7_5 .LUT_INIT=16'b0010110000100100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_26_LC_2_7_5  (
            .in0(N__8725),
            .in1(N__8653),
            .in2(N__8577),
            .in3(N__8773),
            .lcout(\uu2.mem0.w_data_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNIOJJI1_2_LC_2_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNIOJJI1_2_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNIOJJI1_2_LC_2_7_6 .LUT_INIT=16'b1011111110001000;
    LogicCell40 \Lab_UT.dspStr.cnt_RNIOJJI1_2_LC_2_7_6  (
            .in0(N__8563),
            .in1(N__8722),
            .in2(N__10155),
            .in3(N__8657),
            .lcout(Lab_UT_L3_tx_data_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNIPKJI1_2_LC_2_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNIPKJI1_2_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNIPKJI1_2_LC_2_7_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dspStr.cnt_RNIPKJI1_2_LC_2_7_7  (
            .in0(N__8721),
            .in1(N__8652),
            .in2(N__10224),
            .in3(N__8564),
            .lcout(L3_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNILGJI1_2_LC_2_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNILGJI1_2_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNILGJI1_2_LC_2_8_0 .LUT_INIT=16'b1010101010001111;
    LogicCell40 \Lab_UT.dspStr.cnt_RNILGJI1_2_LC_2_8_0  (
            .in0(N__8650),
            .in1(N__8808),
            .in2(N__8745),
            .in3(N__8569),
            .lcout(L3_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIG1C8B_2_LC_2_8_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIG1C8B_2_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIG1C8B_2_LC_2_8_1 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uu2.w_addr_user_RNIG1C8B_2_LC_2_8_1  (
            .in0(N__6968),
            .in1(N__7206),
            .in2(N__7053),
            .in3(N__6897),
            .lcout(\uu2.un27_w_addr_user_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.rdy_LC_2_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.rdy_LC_2_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.rdy_LC_2_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dspStr.rdy_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6933),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13522),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_5_1_LC_2_8_3 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_5_1_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_5_1_LC_2_8_3 .LUT_INIT=16'b0100000000110011;
    LogicCell40 \uu2.un1_w_user_cr_5_1_LC_2_8_3  (
            .in0(N__10197),
            .in1(N__8737),
            .in2(N__8815),
            .in3(N__8649),
            .lcout(\uu2.un1_w_user_cr_5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_3_LC_2_8_4 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_3_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_3_LC_2_8_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uu2.un1_w_user_lf_3_LC_2_8_4  (
            .in0(N__8651),
            .in1(N__8754),
            .in2(N__10163),
            .in3(N__6915),
            .lcout(\uu2.un1_w_user_lfZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_2_LC_2_8_5 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_2_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_2_LC_2_8_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uu2.un1_w_user_cr_2_LC_2_8_5  (
            .in0(N__7037),
            .in1(N__6878),
            .in2(_gnd_net_),
            .in3(N__6903),
            .lcout(\uu2.un1_w_user_crZ0Z_2 ),
            .ltout(\uu2.un1_w_user_crZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un19_w_addr_user_0_LC_2_8_6 .C_ON=1'b0;
    defparam \uu2.un19_w_addr_user_0_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.un19_w_addr_user_0_LC_2_8_6 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \uu2.un19_w_addr_user_0_LC_2_8_6  (
            .in0(N__6891),
            .in1(N__7052),
            .in2(N__6885),
            .in3(N__6967),
            .lcout(\uu2.un19_w_addr_userZ0Z_0 ),
            .ltout(\uu2.un19_w_addr_userZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_2_8_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_2_8_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_15_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6882),
            .in3(N__6879),
            .lcout(\uu2.mem0.w_data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNIIDJI1_2_LC_2_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNIIDJI1_2_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNIIDJI1_2_LC_2_9_0 .LUT_INIT=16'b1111111110110011;
    LogicCell40 \Lab_UT.dspStr.cnt_RNIIDJI1_2_LC_2_9_0  (
            .in0(N__8729),
            .in1(N__8655),
            .in2(N__10369),
            .in3(N__8566),
            .lcout(Lab_UT_L3_tx_data_2_0),
            .ltout(Lab_UT_L3_tx_data_2_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_5_LC_2_9_1 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_5_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_5_LC_2_9_1 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \uu2.un1_w_user_cr_5_LC_2_9_1  (
            .in0(N__8567),
            .in1(N__7062),
            .in2(N__7056),
            .in3(N__8658),
            .lcout(\uu2.un1_w_user_crZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_2_9_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_2_9_2 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_2_9_2  (
            .in0(N__7041),
            .in1(N__8927),
            .in2(_gnd_net_),
            .in3(N__12425),
            .lcout(\uu2.mem0.w_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_2_9_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_2_9_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__12420),
            .in2(N__7020),
            .in3(N__12576),
            .lcout(\uu2.mem0.w_addr_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_2_9_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_2_9_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_21_LC_2_9_4  (
            .in0(N__8731),
            .in1(N__6987),
            .in2(_gnd_net_),
            .in3(N__8656),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_2_9_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_2_9_5 .LUT_INIT=16'b0101000110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_22_LC_2_9_5  (
            .in0(N__8568),
            .in1(N__8730),
            .in2(N__8859),
            .in3(N__8659),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_2_9_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_2_9_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_2_9_6  (
            .in0(N__7130),
            .in1(_gnd_net_),
            .in2(N__12462),
            .in3(N__14998),
            .lcout(\uu2.mem0.w_addr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_2_9_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_2_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(N__12424),
            .in2(_gnd_net_),
            .in3(N__6972),
            .lcout(\uu2.mem0.w_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_3_LC_2_10_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_3_LC_2_10_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_3_LC_2_10_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uu2.w_addr_user_3_LC_2_10_1  (
            .in0(N__8988),
            .in1(_gnd_net_),
            .in2(N__7143),
            .in3(N__7191),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_3C_net ),
            .ce(),
            .sr(N__7164));
    defparam \uu2.w_addr_user_1_LC_2_10_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_1_LC_2_10_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.w_addr_user_1_LC_2_10_2  (
            .in0(N__7190),
            .in1(_gnd_net_),
            .in2(N__8095),
            .in3(N__7133),
            .lcout(\uu2.w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_3C_net ),
            .ce(),
            .sr(N__7164));
    defparam \uu2.w_addr_user_RNIDD1A_5_LC_2_10_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIDD1A_5_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIDD1A_5_LC_2_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_RNIDD1A_5_LC_2_10_3  (
            .in0(N__8987),
            .in1(N__7129),
            .in2(N__9323),
            .in3(N__8082),
            .lcout(),
            .ltout(\uu2.un2_w_addr_user_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIDMJM_2_LC_2_10_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIDMJM_2_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIDMJM_2_LC_2_10_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uu2.w_addr_user_RNIDMJM_2_LC_2_10_4  (
            .in0(N__9365),
            .in1(N__9035),
            .in2(N__7215),
            .in3(N__7212),
            .lcout(\uu2.un2_w_addr_user ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_0_LC_2_10_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_0_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_0_LC_2_10_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_user_0_LC_2_10_5  (
            .in0(_gnd_net_),
            .in1(N__8083),
            .in2(_gnd_net_),
            .in3(N__7189),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_3C_net ),
            .ce(),
            .sr(N__7164));
    defparam \uu2.w_addr_user_2_LC_2_10_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_2_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_2_LC_2_10_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_user_2_LC_2_10_6  (
            .in0(N__7192),
            .in1(N__9036),
            .in2(N__8096),
            .in3(N__7134),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_3C_net ),
            .ce(),
            .sr(N__7164));
    defparam \uu2.w_addr_user_5_LC_2_10_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_5_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_5_LC_2_10_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_user_5_LC_2_10_7  (
            .in0(N__9318),
            .in1(N__9366),
            .in2(N__7101),
            .in3(N__7193),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_3C_net ),
            .ce(),
            .sr(N__7164));
    defparam \uu2.vbuf_w_addr_user.result_1_3_LC_2_11_0 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.result_1_3_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.result_1_3_LC_2_11_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.vbuf_w_addr_user.result_1_3_LC_2_11_0  (
            .in0(N__8094),
            .in1(N__8990),
            .in2(N__9047),
            .in3(N__7132),
            .lcout(\uu2.o_adder_vbuf_w_addr_user_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un425_ci_LC_2_11_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un425_ci_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un425_ci_LC_2_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_4__un425_ci_LC_2_11_7  (
            .in0(N__8989),
            .in1(N__7131),
            .in2(N__9046),
            .in3(N__8093),
            .lcout(\uu2.un425_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_esr_3_LC_2_12_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_3_LC_2_12_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_3_LC_2_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_3_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7071),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13496),
            .ce(N__11352),
            .sr(N__15878));
    defparam \Lab_UT.secuu0.l_count_17_LC_4_4_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_17_LC_4_4_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_17_LC_4_4_1 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \Lab_UT.secuu0.l_count_17_LC_4_4_1  (
            .in0(N__7258),
            .in1(N__7673),
            .in2(N__7311),
            .in3(N__7288),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13535),
            .ce(N__7587),
            .sr(N__15902));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_11__un186_ci_0_LC_4_4_2 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_11__un186_ci_0_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_11__un186_ci_0_LC_4_4_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_11__un186_ci_0_LC_4_4_2  (
            .in0(N__7521),
            .in1(N__7483),
            .in2(_gnd_net_),
            .in3(N__7452),
            .lcout(),
            .ltout(\Lab_UT.secuu0.un186_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_11_LC_4_4_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_11_LC_4_4_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_11_LC_4_4_3 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \Lab_UT.secuu0.l_count_11_LC_4_4_3  (
            .in0(N__7675),
            .in1(N__7367),
            .in2(N__7497),
            .in3(N__11068),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13535),
            .ce(N__7587),
            .sr(N__15902));
    defparam \Lab_UT.secuu0.l_count_16_LC_4_4_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_16_LC_4_4_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_16_LC_4_4_4 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Lab_UT.secuu0.l_count_16_LC_4_4_4  (
            .in0(N__11069),
            .in1(N__7676),
            .in2(N__7290),
            .in3(N__7257),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13535),
            .ce(N__7587),
            .sr(N__15902));
    defparam \Lab_UT.secuu0.l_count_8_LC_4_4_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_8_LC_4_4_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_8_LC_4_4_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.secuu0.l_count_8_LC_4_4_5  (
            .in0(N__7484),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7672),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13535),
            .ce(N__7587),
            .sr(N__15902));
    defparam \Lab_UT.secuu0.l_count_RNIRDS11_3_LC_4_5_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNIRDS11_3_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNIRDS11_3_LC_4_5_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNIRDS11_3_LC_4_5_0  (
            .in0(N__7451),
            .in1(N__7413),
            .in2(N__7310),
            .in3(N__7394),
            .lcout(),
            .ltout(\Lab_UT.secuu0.un4_l_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_RNIOSIV1_18_LC_4_5_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNIOSIV1_18_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNIOSIV1_18_LC_4_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNIOSIV1_18_LC_4_5_1  (
            .in0(N__7226),
            .in1(N__7363),
            .in2(N__7347),
            .in3(N__7344),
            .lcout(\Lab_UT.secuu0.un4_l_count_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_13__un208_ci_0_LC_4_5_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_13__un208_ci_0_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_13__un208_ci_0_LC_4_5_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_13__un208_ci_0_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__7733),
            .in2(_gnd_net_),
            .in3(N__7702),
            .lcout(\Lab_UT.secuu0.un208_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_18__un263_ci_LC_4_5_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_18__un263_ci_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_18__un263_ci_LC_4_5_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_18__un263_ci_LC_4_5_6  (
            .in0(N__7306),
            .in1(N__7289),
            .in2(N__7262),
            .in3(N__7653),
            .lcout(\Lab_UT.secuu0.un263_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_18_LC_4_6_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_18_LC_4_6_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_18_LC_4_6_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \Lab_UT.secuu0.l_count_18_LC_4_6_0  (
            .in0(N__7233),
            .in1(N__7227),
            .in2(_gnd_net_),
            .in3(N__11072),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13523),
            .ce(N__7585),
            .sr(N__15900));
    defparam \Lab_UT.secuu0.l_count_12_LC_4_6_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_12_LC_4_6_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_12_LC_4_6_4 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \Lab_UT.secuu0.l_count_12_LC_4_6_4  (
            .in0(N__7682),
            .in1(N__7703),
            .in2(N__7737),
            .in3(N__11070),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13523),
            .ce(N__7585),
            .sr(N__15900));
    defparam \Lab_UT.secuu0.l_count_13_LC_4_6_7 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_13_LC_4_6_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_13_LC_4_6_7 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \Lab_UT.secuu0.l_count_13_LC_4_6_7  (
            .in0(N__11071),
            .in1(N__7683),
            .in2(N__7605),
            .in3(N__7611),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13523),
            .ce(N__7585),
            .sr(N__15900));
    defparam \Lab_UT.secuu0.l_precount_0_LC_4_7_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_precount_0_LC_4_7_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_precount_0_LC_4_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.secuu0.l_precount_0_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7540),
            .lcout(\Lab_UT.secuu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13516),
            .ce(),
            .sr(N__15877));
    defparam \uu2.r_addr_5_LC_4_7_2 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_4_7_2 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_5_LC_4_7_2  (
            .in0(N__7848),
            .in1(N__7940),
            .in2(N__7919),
            .in3(N__11192),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13516),
            .ce(),
            .sr(N__15877));
    defparam \uu2.r_addr_4_LC_4_7_5 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_4_7_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_4_7_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.r_addr_4_LC_4_7_5  (
            .in0(N__11191),
            .in1(N__7847),
            .in2(_gnd_net_),
            .in3(N__7914),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13516),
            .ce(),
            .sr(N__15877));
    defparam \uu2.r_addr_0_LC_4_7_6 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_4_7_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_4_7_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.r_addr_0_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(N__11255),
            .in2(_gnd_net_),
            .in3(N__11190),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13516),
            .ce(),
            .sr(N__15877));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un425_ci_LC_4_8_0 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un425_ci_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un425_ci_LC_4_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un425_ci_LC_4_8_0  (
            .in0(N__11104),
            .in1(N__11314),
            .in2(N__7801),
            .in3(N__11253),
            .lcout(\uu2.un425_ci_0 ),
            .ltout(\uu2.un425_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_6_LC_4_8_1 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_4_8_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.r_addr_esr_6_LC_4_8_1  (
            .in0(N__7939),
            .in1(N__7918),
            .in2(N__7524),
            .in3(N__7871),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13510),
            .ce(N__11341),
            .sr(N__15874));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un469_ci_0_LC_4_8_2 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un469_ci_0_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un469_ci_0_LC_4_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un469_ci_0_LC_4_8_2  (
            .in0(_gnd_net_),
            .in1(N__7822),
            .in2(_gnd_net_),
            .in3(N__7869),
            .lcout(),
            .ltout(\uu2.vbuf_raddr.un469_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_8_LC_4_8_3 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_4_8_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_4_8_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_8_LC_4_8_3  (
            .in0(N__7961),
            .in1(N__7884),
            .in2(N__7971),
            .in3(N__7845),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13510),
            .ce(N__11341),
            .sr(N__15874));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un447_ci_3_LC_4_8_4 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un447_ci_3_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un447_ci_3_LC_4_8_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un447_ci_3_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(N__7938),
            .in2(_gnd_net_),
            .in3(N__7904),
            .lcout(\uu2.vbuf_raddr.un447_ci_3 ),
            .ltout(\uu2.vbuf_raddr.un447_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_7_LC_4_8_5 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_4_8_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_7_LC_4_8_5  (
            .in0(N__7870),
            .in1(N__7823),
            .in2(N__7851),
            .in3(N__7846),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13510),
            .ce(N__11341),
            .sr(N__15874));
    defparam \uu2.r_addr_esr_3_LC_4_8_6 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_4_8_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_4_8_6  (
            .in0(N__11105),
            .in1(N__11315),
            .in2(N__7802),
            .in3(N__11254),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13510),
            .ce(N__11341),
            .sr(N__15874));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_9_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_4_9_0  (
            .in0(N__12476),
            .in1(N__7779),
            .in2(_gnd_net_),
            .in3(N__7746),
            .lcout(\uu2.mem0.w_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_9_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_9_1 .LUT_INIT=16'b1010101000000011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_4_9_1  (
            .in0(N__7764),
            .in1(N__9235),
            .in2(N__8931),
            .in3(N__12478),
            .lcout(\uu2.mem0.w_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_4_9_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_4_9_2 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_17_LC_4_9_2  (
            .in0(N__8918),
            .in1(_gnd_net_),
            .in2(N__9236),
            .in3(N__16202),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_4_9_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_4_9_3 .LUT_INIT=16'b0001000000110011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_37_LC_4_9_3  (
            .in0(N__11439),
            .in1(N__12475),
            .in2(N__7989),
            .in3(N__8181),
            .lcout(),
            .ltout(\uu2.mem0.G_14_0_a6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_4_9_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_4_9_4 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_24_LC_4_9_4  (
            .in0(N__10419),
            .in1(N__10560),
            .in2(N__7740),
            .in3(N__9096),
            .lcout(),
            .ltout(\uu2.mem0.N_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_9_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_9_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_4_9_5  (
            .in0(N__11748),
            .in1(N__8940),
            .in2(N__8016),
            .in3(N__9249),
            .lcout(\uu2.mem0.w_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_4_9_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_4_9_6 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_18_LC_4_9_6  (
            .in0(N__8919),
            .in1(_gnd_net_),
            .in2(N__9237),
            .in3(N__16203),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_9_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_9_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(N__8007),
            .in2(N__7998),
            .in3(N__12477),
            .lcout(\uu2.mem0.w_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNII1IB1_5_LC_4_10_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNII1IB1_5_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNII1IB1_5_LC_4_10_0 .LUT_INIT=16'b0001001000010000;
    LogicCell40 \uu2.w_addr_displaying_RNII1IB1_5_LC_4_10_0  (
            .in0(N__12229),
            .in1(N__12562),
            .in2(N__12322),
            .in3(N__16287),
            .lcout(\uu2.bitmap_pmux_1_1_a8_1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_4_10_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_4_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_49_LC_4_10_1  (
            .in0(N__16288),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12563),
            .lcout(\uu2.mem0.G_14_0_a6_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_10_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_10_2 .LUT_INIT=16'b0101110101011111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_4_10_2  (
            .in0(N__8151),
            .in1(N__9135),
            .in2(N__12482),
            .in3(N__9108),
            .lcout(\uu2.mem0.w_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI979P_3_LC_4_10_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI979P_3_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI979P_3_LC_4_10_3 .LUT_INIT=16'b1101111111111011;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI979P_3_LC_4_10_3  (
            .in0(N__13083),
            .in1(N__14832),
            .in2(N__14987),
            .in3(N__14313),
            .lcout(\uu2.N_326_0 ),
            .ltout(\uu2.N_326_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0QUP1_6_LC_4_10_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0QUP1_6_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0QUP1_6_LC_4_10_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \uu2.w_addr_displaying_RNI0QUP1_6_LC_4_10_4  (
            .in0(N__12230),
            .in1(N__12561),
            .in2(N__7974),
            .in3(N__16286),
            .lcout(\uu2.bitmap_pmux_1_1_a8_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI28SI1_7_LC_4_10_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI28SI1_7_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI28SI1_7_LC_4_10_5 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI28SI1_7_LC_4_10_5  (
            .in0(N__13856),
            .in1(N__14010),
            .in2(N__13035),
            .in3(N__14253),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_1_1_a8_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNITAMH5_7_LC_4_10_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNITAMH5_7_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNITAMH5_7_LC_4_10_6 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \uu2.w_addr_displaying_fast_RNITAMH5_7_LC_4_10_6  (
            .in0(N__8202),
            .in1(N__8196),
            .in2(N__8190),
            .in3(N__8187),
            .lcout(\uu2.bitmap_pmux_1_1_1_tz ),
            .ltout(\uu2.bitmap_pmux_1_1_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_4_10_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_4_10_7 .LUT_INIT=16'b1111000010010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_29_LC_4_10_7  (
            .in0(N__16289),
            .in1(N__12564),
            .in2(N__8175),
            .in3(N__11435),
            .lcout(\uu2.mem0.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_4_11_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_4_11_0 .LUT_INIT=16'b0000111100010001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_25_LC_4_11_0  (
            .in0(N__9217),
            .in1(N__8926),
            .in2(N__8172),
            .in3(N__12466),
            .lcout(\uu2.mem0.w_data_1_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_wr_en_0_i_LC_4_11_2 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_4_11_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_4_11_2  (
            .in0(N__8141),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12467),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_4_11_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_4_11_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_4_11_3  (
            .in0(N__12468),
            .in1(N__8100),
            .in2(_gnd_net_),
            .in3(N__16200),
            .lcout(\uu2.mem0.w_addr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_LC_4_11_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_LC_4_11_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_LC_4_11_7 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.w_addr_displaying_1_LC_4_11_7  (
            .in0(N__16098),
            .in1(N__16201),
            .in2(_gnd_net_),
            .in3(N__14961),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1C_net ),
            .ce(),
            .sr(N__15848));
    defparam \uu2.r_data_reg_esr_1_LC_4_12_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_1_LC_4_12_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_1_LC_4_12_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uu2.r_data_reg_esr_1_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__8046),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13489),
            .ce(N__11348),
            .sr(N__15881));
    defparam \uu2.r_data_reg_esr_2_LC_4_12_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_2_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_2_LC_4_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_2_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8037),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13489),
            .ce(N__11348),
            .sr(N__15881));
    defparam \uu2.r_data_reg_esr_0_LC_4_12_3 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_0_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_0_LC_4_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_0_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8028),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13489),
            .ce(N__11348),
            .sr(N__15881));
    defparam \uu2.r_data_reg_esr_4_LC_4_12_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_4_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_4_LC_4_12_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uu2.r_data_reg_esr_4_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__8289),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13489),
            .ce(N__11348),
            .sr(N__15881));
    defparam \uu2.r_data_reg_esr_5_LC_4_12_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_5_LC_4_12_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_5_LC_4_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_5_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8280),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13489),
            .ce(N__11348),
            .sr(N__15881));
    defparam \uu2.r_data_reg_esr_6_LC_4_12_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_6_LC_4_12_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_6_LC_4_12_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_esr_6_LC_4_12_6  (
            .in0(N__8271),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13489),
            .ce(N__11348),
            .sr(N__15881));
    defparam \uu2.r_data_reg_esr_7_LC_4_12_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_7_LC_4_12_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_7_LC_4_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_esr_7_LC_4_12_7  (
            .in0(N__8262),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13489),
            .ce(N__11348),
            .sr(N__15881));
    defparam \buart.Z_tx.shifter_1_LC_4_13_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_4_13_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_1_LC_4_13_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \buart.Z_tx.shifter_1_LC_4_13_0  (
            .in0(N__11223),
            .in1(_gnd_net_),
            .in2(N__8253),
            .in3(N__8214),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13486),
            .ce(N__9570),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_0_LC_4_13_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_0_LC_4_13_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_tx.shifter_0_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__8244),
            .in2(_gnd_net_),
            .in3(N__11221),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13486),
            .ce(N__9570),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.uart_tx_LC_4_13_2 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.uart_tx_LC_4_13_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \buart.Z_tx.uart_tx_LC_4_13_2  (
            .in0(N__11222),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8238),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13486),
            .ce(N__9570),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_2_LC_4_13_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_4_13_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_2_LC_4_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \buart.Z_tx.shifter_2_LC_4_13_3  (
            .in0(N__8220),
            .in1(N__8346),
            .in2(_gnd_net_),
            .in3(N__11224),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13486),
            .ce(N__9570),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_3_LC_4_13_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_4_13_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_3_LC_4_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \buart.Z_tx.shifter_3_LC_4_13_4  (
            .in0(N__11225),
            .in1(N__8208),
            .in2(_gnd_net_),
            .in3(N__8328),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13486),
            .ce(N__9570),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_4_LC_4_13_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_4_LC_4_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \buart.Z_tx.shifter_4_LC_4_13_5  (
            .in0(N__8340),
            .in1(N__8316),
            .in2(_gnd_net_),
            .in3(N__11226),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13486),
            .ce(N__9570),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_5_LC_4_13_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_4_13_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_5_LC_4_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \buart.Z_tx.shifter_5_LC_4_13_6  (
            .in0(N__11227),
            .in1(N__8322),
            .in2(_gnd_net_),
            .in3(N__8304),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13486),
            .ce(N__9570),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_6_LC_4_13_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_4_13_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_6_LC_4_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \buart.Z_tx.shifter_6_LC_4_13_7  (
            .in0(N__9159),
            .in1(N__8310),
            .in2(_gnd_net_),
            .in3(N__11228),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13486),
            .ce(N__9570),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_2_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_2_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_2_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_5_3_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_5_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__10105),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_5_3_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_5_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_5_3_1  (
            .in0(_gnd_net_),
            .in1(N__8405),
            .in2(_gnd_net_),
            .in3(N__8298),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_5_3_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_5_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_5_3_2  (
            .in0(_gnd_net_),
            .in1(N__10069),
            .in2(_gnd_net_),
            .in3(N__8295),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_5_3_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_5_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__10013),
            .in2(_gnd_net_),
            .in3(N__8292),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_4_LC_5_3_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_4_LC_5_3_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_e_0_4_LC_5_3_4 .LUT_INIT=16'b0001101101001110;
    LogicCell40 \buart.Z_rx.bitcount_e_0_4_LC_5_3_4  (
            .in0(N__8885),
            .in1(N__8427),
            .in2(N__9897),
            .in3(N__8433),
            .lcout(buart__rx_bitcount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13536),
            .ce(N__9825),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNI2B26_4_LC_5_4_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNI2B26_4_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNI2B26_4_LC_5_4_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNI2B26_4_LC_5_4_0  (
            .in0(N__8404),
            .in1(N__10070),
            .in2(N__10023),
            .in3(N__8426),
            .lcout(),
            .ltout(\buart.Z_rx.N_144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNIBJOC_0_LC_5_4_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNIBJOC_0_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNIBJOC_0_LC_5_4_1 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNIBJOC_0_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(N__9930),
            .in2(N__8430),
            .in3(N__10111),
            .lcout(\buart.Z_rx.N_41_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_i_0_o2_4_LC_5_4_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_i_0_o2_4_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_2_i_0_o2_4_LC_5_4_3 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \resetGen.reset_count_2_i_0_o2_4_LC_5_4_3  (
            .in0(N__8425),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8403),
            .lcout(N_118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_1_LC_5_4_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_1_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_e_0_1_LC_5_4_4 .LUT_INIT=16'b0001101101001110;
    LogicCell40 \buart.Z_rx.bitcount_e_0_1_LC_5_4_4  (
            .in0(N__8880),
            .in1(N__8412),
            .in2(N__9888),
            .in3(N__8406),
            .lcout(buart__rx_bitcount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13529),
            .ce(N__9824),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_2_LC_5_4_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_2_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_e_0_2_LC_5_4_5 .LUT_INIT=16'b0011001101011010;
    LogicCell40 \buart.Z_rx.bitcount_e_0_2_LC_5_4_5  (
            .in0(N__10071),
            .in1(N__9875),
            .in2(N__8385),
            .in3(N__8881),
            .lcout(buart__rx_bitcount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13529),
            .ce(N__9824),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_3_LC_5_4_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_3_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_e_0_3_LC_5_4_6 .LUT_INIT=16'b0101001101011100;
    LogicCell40 \buart.Z_rx.bitcount_e_0_3_LC_5_4_6  (
            .in0(N__9873),
            .in1(N__8376),
            .in2(N__8886),
            .in3(N__10014),
            .lcout(buart__rx_bitcount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13529),
            .ce(N__9824),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_0_LC_5_4_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_0_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_e_0_0_LC_5_4_7 .LUT_INIT=16'b0011001101011010;
    LogicCell40 \buart.Z_rx.bitcount_e_0_0_LC_5_4_7  (
            .in0(N__10112),
            .in1(N__9874),
            .in2(N__8369),
            .in3(N__8879),
            .lcout(buart__rx_bitcount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13529),
            .ce(N__9824),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_4_LC_5_5_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_4_LC_5_5_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_4_LC_5_5_0  (
            .in0(N__8492),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13524),
            .ce(N__13570),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_i_0_a3_5_4_LC_5_5_2 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_i_0_a3_5_4_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_2_i_0_a3_5_4_LC_5_5_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \resetGen.reset_count_2_i_0_a3_5_4_LC_5_5_2  (
            .in0(N__8491),
            .in1(N__9658),
            .in2(N__9686),
            .in3(N__13592),
            .lcout(),
            .ltout(\resetGen.reset_count_2_i_0_a3_5Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_i_0_a3_4_LC_5_5_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_i_0_a3_4_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_2_i_0_a3_4_LC_5_5_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \resetGen.reset_count_2_i_0_a3_4_LC_5_5_3  (
            .in0(N__8478),
            .in1(N__8472),
            .in2(N__8502),
            .in3(N__9969),
            .lcout(\resetGen.N_133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_5_LC_5_5_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_5_LC_5_5_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_5_LC_5_5_4  (
            .in0(N__9682),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13524),
            .ce(N__13570),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_7_LC_5_5_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_7_LC_5_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8466),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13524),
            .ce(N__13570),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_i_0_a3_6_4_LC_5_5_7 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_i_0_a3_6_4_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_2_i_0_a3_6_4_LC_5_5_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \resetGen.reset_count_2_i_0_a3_6_4_LC_5_5_7  (
            .in0(N__13615),
            .in1(N__10009),
            .in2(N__9614),
            .in3(N__10063),
            .lcout(\resetGen.reset_count_2_i_0_a3_6Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_i_0_a3_4_4_LC_5_6_2 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_i_0_a3_4_4_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_2_i_0_a3_4_4_LC_5_6_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \resetGen.reset_count_2_i_0_a3_4_4_LC_5_6_2  (
            .in0(N__10114),
            .in1(N__9713),
            .in2(_gnd_net_),
            .in3(N__9634),
            .lcout(\resetGen.reset_count_2_i_0_a3_4Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_1_LC_5_6_3 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.hh_1_LC_5_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8451),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13517),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_LC_5_6_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_LC_5_6_4 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNI8RI7_0_LC_5_6_4  (
            .in0(N__10113),
            .in1(N__10072),
            .in2(N__10030),
            .in3(N__9970),
            .lcout(\buart.Z_rx.N_129 ),
            .ltout(\buart.Z_rx.N_129_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_RNIVHME_0_LC_5_6_5 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNIVHME_0_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNIVHME_0_LC_5_6_5 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \buart.Z_rx.hh_RNIVHME_0_LC_5_6_5  (
            .in0(_gnd_net_),
            .in1(N__8465),
            .in2(N__8454),
            .in3(N__8450),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.Lab3U00.q_esr_ctle_7_LC_5_6_6 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_ctle_7_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.Lab3U00.q_esr_ctle_7_LC_5_6_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_ctle_7_LC_5_6_6  (
            .in0(N__9945),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15917),
            .lcout(\Lab_UT.Lab3U00.bu_rx_data_rdy_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNIGM5F_0_LC_5_6_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNIGM5F_0_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNIGM5F_0_LC_5_6_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNIGM5F_0_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__9944),
            .in2(_gnd_net_),
            .in3(N__9911),
            .lcout(\buart.Z_rx.N_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec1.segmentUQ_0_LC_5_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dec1.segmentUQ_0_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec1.segmentUQ_0_LC_5_7_0 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \Lab_UT.dec1.segmentUQ_0_LC_5_7_0  (
            .in0(N__14198),
            .in1(N__17335),
            .in2(N__14120),
            .in3(N__15646),
            .lcout(L3_segment2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_3_LC_5_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_3_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_3_LC_5_7_2 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \Lab_UT.dictrluu0.dicfsm.cState_RNO_3_LC_5_7_2  (
            .in0(N__8858),
            .in1(N__10364),
            .in2(N__8820),
            .in3(N__10316),
            .lcout(\Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dek.det_N_0_a3_1_LC_5_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dek.det_N_0_a3_1_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrluu0.dek.det_N_0_a3_1_LC_5_7_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.dictrluu0.dek.det_N_0_a3_1_LC_5_7_4  (
            .in0(N__8857),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8816),
            .lcout(\Lab_UT.dictrluu0.N_103_1 ),
            .ltout(\Lab_UT.dictrluu0.N_103_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_1_LC_5_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_1_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_1_LC_5_7_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrluu0.dicfsm.cState_RNO_1_LC_5_7_5  (
            .in0(N__10365),
            .in1(N__10312),
            .in2(N__8784),
            .in3(N__8781),
            .lcout(\Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec3.g0_0_LC_5_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dec3.g0_0_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec3.g0_0_LC_5_7_7 .LUT_INIT=16'b0110000100000010;
    LogicCell40 \Lab_UT.dec3.g0_0_LC_5_7_7  (
            .in0(N__15187),
            .in1(N__17061),
            .in2(N__15102),
            .in3(N__17450),
            .lcout(N_52_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_3_1_LC_5_8_0 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_3_1_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_3_1_LC_5_8_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uu2.un1_w_user_lf_3_1_LC_5_8_0  (
            .in0(N__10182),
            .in1(N__8743),
            .in2(_gnd_net_),
            .in3(N__8575),
            .lcout(\uu2.un1_w_user_lf_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_5_8_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_5_8_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_44_LC_5_8_1  (
            .in0(N__8744),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10183),
            .lcout(),
            .ltout(\uu2.mem0.N_26_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_5_8_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_5_8_2 .LUT_INIT=16'b0010001000001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_31_LC_5_8_2  (
            .in0(N__12427),
            .in1(N__8667),
            .in2(N__8580),
            .in3(N__8576),
            .lcout(\uu2.mem0.G_14_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.Lab3U00.q_esr_1_LC_5_8_3 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_1_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_1_LC_5_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_1_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13626),
            .lcout(Lab_UT_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13501),
            .ce(N__9082),
            .sr(N__15876));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_5_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_5_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_5_8_4  (
            .in0(N__12428),
            .in1(N__9048),
            .in2(_gnd_net_),
            .in3(N__11703),
            .lcout(\uu2.mem0.w_addr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI80631_4_LC_5_8_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI80631_4_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI80631_4_LC_5_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI80631_4_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(N__13995),
            .in2(_gnd_net_),
            .in3(N__13002),
            .lcout(\uu2.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_5_8_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_5_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_5_8_7  (
            .in0(N__12840),
            .in1(N__8994),
            .in2(_gnd_net_),
            .in3(N__12429),
            .lcout(\uu2.mem0.w_addr_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec1.g0_i_LC_5_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dec1.g0_i_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec1.g0_i_LC_5_9_0 .LUT_INIT=16'b1001111011111011;
    LogicCell40 \Lab_UT.dec1.g0_i_LC_5_9_0  (
            .in0(N__17342),
            .in1(N__14199),
            .in2(N__14121),
            .in3(N__15653),
            .lcout(L3_segment2_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_5_9_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_5_9_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_32_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__8917),
            .in2(_gnd_net_),
            .in3(N__16183),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_32_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_5_9_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_5_9_3 .LUT_INIT=16'b1100110011111110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_19_LC_5_9_3  (
            .in0(N__9228),
            .in1(N__8949),
            .in2(N__8943),
            .in3(N__12471),
            .lcout(\uu2.mem0.G_14_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI6NLE_7_LC_5_9_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI6NLE_7_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI6NLE_7_LC_5_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI6NLE_7_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(N__13847),
            .in2(_gnd_net_),
            .in3(N__14246),
            .lcout(),
            .ltout(\uu2.N_329_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIV60G2_2_LC_5_9_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIV60G2_2_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIV60G2_2_LC_5_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIV60G2_2_LC_5_9_5  (
            .in0(N__10377),
            .in1(N__11698),
            .in2(N__8934),
            .in3(N__14988),
            .lcout(\uu2.Z_decfrac105_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_5_9_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_5_9_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_57_LC_5_9_6  (
            .in0(N__13791),
            .in1(N__9153),
            .in2(_gnd_net_),
            .in3(N__9144),
            .lcout(),
            .ltout(\uu2.mem0.N_2159_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_5_9_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_5_9_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_50_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(N__14340),
            .in2(N__9138),
            .in3(N__13665),
            .lcout(\uu2.mem0.N_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_5_10_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_5_10_0 .LUT_INIT=16'b0010101000001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_20_LC_5_10_0  (
            .in0(N__11715),
            .in1(N__9243),
            .in2(N__9195),
            .in3(N__10414),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI0OT22_4_LC_5_10_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI0OT22_4_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI0OT22_4_LC_5_10_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI0OT22_4_LC_5_10_1  (
            .in0(N__9180),
            .in1(N__9129),
            .in2(_gnd_net_),
            .in3(N__12657),
            .lcout(\uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4 ),
            .ltout(\uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_5_10_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_5_10_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_41_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__9186),
            .in2(N__9120),
            .in3(N__14425),
            .lcout(\uu2.mem0.un1_segment3_m2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_5_10_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_5_10_3 .LUT_INIT=16'b0111011101110111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_28_LC_5_10_3  (
            .in0(N__11597),
            .in1(N__10547),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\uu2.mem0.N_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_5_10_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_5_10_4 .LUT_INIT=16'b1110110011101111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_16_LC_5_10_4  (
            .in0(N__10500),
            .in1(N__9117),
            .in2(N__9111),
            .in3(N__10413),
            .lcout(\uu2.mem0.bitmap_pmux_1_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_5_10_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_5_10_5 .LUT_INIT=16'b1111101100000001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_38_LC_5_10_5  (
            .in0(N__11596),
            .in1(N__12732),
            .in2(N__12645),
            .in3(N__9102),
            .lcout(\uu2.mem0.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_5_10_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_5_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_46_LC_5_10_6  (
            .in0(N__9267),
            .in1(N__14426),
            .in2(_gnd_net_),
            .in3(N__10526),
            .lcout(\uu2.mem0.un1_segment3_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_5_10_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_5_10_7 .LUT_INIT=16'b1000000011110111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_27_LC_5_10_7  (
            .in0(N__10548),
            .in1(N__11598),
            .in2(N__10418),
            .in3(N__10386),
            .lcout(\uu2.mem0.un1_segment3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_5_11_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_5_11_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_34_LC_5_11_0  (
            .in0(N__11589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10546),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIHKAF2_0_8_LC_5_11_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIHKAF2_0_8_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIHKAF2_0_8_LC_5_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIHKAF2_0_8_LC_5_11_1  (
            .in0(N__15366),
            .in1(N__12565),
            .in2(N__9279),
            .in3(N__12819),
            .lcout(\uu2.Z_decfrac106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_5_11_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_5_11_3 .LUT_INIT=16'b1011101111111010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_47_LC_5_11_3  (
            .in0(N__12644),
            .in1(N__14400),
            .in2(N__12728),
            .in3(N__11588),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_47_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_5_11_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_5_11_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_35_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__9204),
            .in2(N__9198),
            .in3(N__9171),
            .lcout(\uu2.mem0.un1_segment3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_5_11_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_5_11_5 .LUT_INIT=16'b1101111101111001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_55_LC_5_11_5  (
            .in0(N__16682),
            .in1(N__16966),
            .in2(N__16784),
            .in3(N__16875),
            .lcout(\uu2.mem0.N_2160_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec3.segmentUQ_i_0_LC_5_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dec3.segmentUQ_i_0_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec3.segmentUQ_i_0_LC_5_11_6 .LUT_INIT=16'b0100100100010000;
    LogicCell40 \Lab_UT.dec3.segmentUQ_i_0_LC_5_11_6  (
            .in0(N__17064),
            .in1(N__15095),
            .in2(N__15189),
            .in3(N__17449),
            .lcout(N_52),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_5_11_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_5_11_7 .LUT_INIT=16'b0001000101010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_48_LC_5_11_7  (
            .in0(N__12643),
            .in1(N__14399),
            .in2(N__12727),
            .in3(N__11587),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_7_LC_5_12_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_7_LC_5_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \buart.Z_tx.shifter_7_LC_5_12_0  (
            .in0(N__11234),
            .in1(N__9165),
            .in2(_gnd_net_),
            .in3(N__9384),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13487),
            .ce(N__9560),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_8_LC_5_12_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_8_LC_5_12_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \buart.Z_tx.shifter_8_LC_5_12_1  (
            .in0(N__9390),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11233),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13487),
            .ce(N__9560),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_5_12_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_5_12_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_5_12_2  (
            .in0(N__12470),
            .in1(_gnd_net_),
            .in2(N__9378),
            .in3(N__13782),
            .lcout(\uu2.mem0.w_addr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_5_12_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_5_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_5_12_4  (
            .in0(N__12469),
            .in1(N__9327),
            .in2(_gnd_net_),
            .in3(N__12293),
            .lcout(\uu2.mem0.w_addr_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI362A1_3_LC_5_12_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI362A1_3_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI362A1_3_LC_5_12_6 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \uu2.w_addr_displaying_RNI362A1_3_LC_5_12_6  (
            .in0(N__15365),
            .in1(N__12796),
            .in2(_gnd_net_),
            .in3(N__14463),
            .lcout(\uu2.w_addr_displaying_RNI362A1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI50L01_0_2_LC_5_13_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI50L01_0_2_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI50L01_0_2_LC_5_13_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uu2.w_addr_displaying_RNI50L01_0_2_LC_5_13_0  (
            .in0(N__11694),
            .in1(N__16193),
            .in2(_gnd_net_),
            .in3(N__14975),
            .lcout(\uu2.Z_decfrac106_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_5_13_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_5_13_6 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_56_LC_5_13_6  (
            .in0(N__16971),
            .in1(N__16874),
            .in2(N__16788),
            .in3(N__16683),
            .lcout(\uu2.mem0.N_2160_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_1_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_1_0  (
            .in0(_gnd_net_),
            .in1(N__9430),
            .in2(N__9411),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_1_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_6_1_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_6_1_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_6_1_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_6_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9462),
            .in3(N__9255),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__13540),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_6_1_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_6_1_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_6_1_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_6_1_2  (
            .in0(N__10672),
            .in1(N__9449),
            .in2(_gnd_net_),
            .in3(N__9252),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__13540),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_6_1_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_6_1_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_6_1_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_6_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9489),
            .in3(N__9510),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__13540),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_6_1_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_6_1_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_6_1_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_6_1_4  (
            .in0(N__10673),
            .in1(_gnd_net_),
            .in2(N__9501),
            .in3(N__9507),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__13540),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_6_1_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_6_1_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_6_1_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_6_1_5  (
            .in0(N__9476),
            .in1(N__10671),
            .in2(_gnd_net_),
            .in3(N__9504),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13540),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_6_1_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_6_1_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_6_1_6  (
            .in0(N__9497),
            .in1(N__9485),
            .in2(N__9477),
            .in3(N__9458),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_6_1_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_6_1_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_6_1_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_6_1_7  (
            .in0(N__9406),
            .in1(N__9429),
            .in2(N__9450),
            .in3(N__9438),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_0_LC_6_2_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_6_2_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_0_LC_6_2_0 .LUT_INIT=16'b0000110100000010;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_6_2_0  (
            .in0(N__10670),
            .in1(N__10812),
            .in2(N__11189),
            .in3(N__10700),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13532),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_6_2_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_6_2_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9431),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13532),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_6_2_2 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_6_2_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_6_2_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_6_2_2  (
            .in0(N__9432),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9410),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13532),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_6_2_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_6_2_3 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_6_2_3  (
            .in0(N__10715),
            .in1(N__10811),
            .in2(_gnd_net_),
            .in3(N__10669),
            .lcout(\buart.Z_tx.un1_bitcount_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_6_3_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_6_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_6_3_0  (
            .in0(_gnd_net_),
            .in1(N__9527),
            .in2(N__9762),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_6_3_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_6_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_6_3_1  (
            .in0(_gnd_net_),
            .in1(N__9732),
            .in2(_gnd_net_),
            .in3(N__9591),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_6_3_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_6_3_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_6_3_2  (
            .in0(N__9889),
            .in1(N__9540),
            .in2(_gnd_net_),
            .in3(N__9588),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__13527),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_6_3_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_6_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_6_3_3  (
            .in0(_gnd_net_),
            .in1(N__9791),
            .in2(_gnd_net_),
            .in3(N__9585),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_6_3_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_6_3_4 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_6_3_4  (
            .in0(N__9777),
            .in1(N__9934),
            .in2(N__9896),
            .in3(N__9582),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13527),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_6_3_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_6_3_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_6_3_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_6_3_6  (
            .in0(N__9792),
            .in1(N__9935),
            .in2(N__9579),
            .in3(N__9879),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13527),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIV5CT5_3_LC_6_4_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIV5CT5_3_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIV5CT5_3_LC_6_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \buart.Z_tx.bitcount_RNIV5CT5_3_LC_6_4_0  (
            .in0(N__10674),
            .in1(N__11922),
            .in2(_gnd_net_),
            .in3(N__10815),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_4_1 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_6_4_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_6_4_1  (
            .in0(N__9760),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9871),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13521),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_6_4_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_6_4_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_6_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_6_4_2  (
            .in0(N__9870),
            .in1(N__9526),
            .in2(_gnd_net_),
            .in3(N__9761),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13521),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_6_4_3 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_6_4_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_6_4_3  (
            .in0(N__9539),
            .in1(N__9730),
            .in2(N__9528),
            .in3(N__9790),
            .lcout(),
            .ltout(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_6_4_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_6_4_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_6_4_4  (
            .in0(_gnd_net_),
            .in1(N__9776),
            .in2(N__9765),
            .in3(N__9759),
            .lcout(\buart.Z_rx.ser_clk ),
            .ltout(\buart.Z_rx.ser_clk_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_6_4_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_6_4_5 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_6_4_5  (
            .in0(N__9741),
            .in1(N__9731),
            .in2(N__9735),
            .in3(N__9872),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13521),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_6_4_7 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_6_4_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_6_4_7 .LUT_INIT=16'b0101000001000001;
    LogicCell40 \resetGen.reset_count_3_LC_6_4_7  (
            .in0(N__10838),
            .in1(N__10881),
            .in2(N__10956),
            .in3(N__10962),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13521),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_6_LC_6_5_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_6_LC_6_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9709),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13513),
            .ce(N__13577),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_LC_6_5_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_1_LC_6_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9659),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13513),
            .ce(N__13577),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_2_LC_6_5_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_6_5_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_2_LC_6_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9610),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13513),
            .ce(N__13577),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_3_LC_6_5_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_6_5_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_3_LC_6_5_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_3_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(N__9635),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13513),
            .ce(N__13577),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dek.det_N_0_o2_LC_6_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dek.det_N_0_o2_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrluu0.dek.det_N_0_o2_LC_6_6_0 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \Lab_UT.dictrluu0.dek.det_N_0_o2_LC_6_6_0  (
            .in0(N__10195),
            .in1(N__10159),
            .in2(N__10128),
            .in3(N__10226),
            .lcout(\Lab_UT.dictrluu0.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_0_LC_6_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_0_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_0_LC_6_6_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrluu0.dicfsm.cState_RNO_0_LC_6_6_1  (
            .in0(N__10227),
            .in1(N__10196),
            .in2(N__10164),
            .in3(N__10127),
            .lcout(\Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.Lab3U01.q_0_LC_6_6_2 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U01.q_0_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U01.q_0_LC_6_6_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.Lab3U01.q_0_LC_6_6_2  (
            .in0(N__10116),
            .in1(N__10074),
            .in2(N__10032),
            .in3(N__9972),
            .lcout(\Lab_UT.rx_data_rdy ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13505),
            .ce(),
            .sr(N__15882));
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_0_LC_6_6_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_0_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_0_LC_6_6_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNI8RI7_0_0_LC_6_6_6  (
            .in0(N__10115),
            .in1(N__10073),
            .in2(N__10031),
            .in3(N__9971),
            .lcout(bu_rx_data_rdy),
            .ltout(bu_rx_data_rdy_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNII0231_0_LC_6_6_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNII0231_0_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNII0231_0_LC_6_6_7 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNII0231_0_LC_6_6_7  (
            .in0(N__9936),
            .in1(N__9912),
            .in2(N__9900),
            .in3(N__9845),
            .lcout(\buart.Z_rx.bitcount_e_0_RNII0231Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec3.segmentUQ_0_6_LC_6_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dec3.segmentUQ_0_6_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec3.segmentUQ_0_6_LC_6_7_1 .LUT_INIT=16'b1111110111101110;
    LogicCell40 \Lab_UT.dec3.segmentUQ_0_6_LC_6_7_1  (
            .in0(N__15131),
            .in1(N__17003),
            .in2(N__17421),
            .in3(N__15047),
            .lcout(),
            .ltout(Lab_UT_dec3_segmentUQ_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment4_1_am_LC_6_7_2 .C_ON=1'b0;
    defparam \uu2.un1_segment4_1_am_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_1_am_LC_6_7_2 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \uu2.un1_segment4_1_am_LC_6_7_2  (
            .in0(N__15049),
            .in1(N__9801),
            .in2(N__9804),
            .in3(N__15133),
            .lcout(\uu2.un1_segment4_1_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpmtens.q_RNIRE5_1_LC_6_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmtens.q_RNIRE5_1_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpmtens.q_RNIRE5_1_LC_6_7_3 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.didpuu0.didpmtens.q_RNIRE5_1_LC_6_7_3  (
            .in0(_gnd_net_),
            .in1(N__17002),
            .in2(_gnd_net_),
            .in3(N__17393),
            .lcout(N_71),
            .ltout(N_71_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpmtens.q_2_LC_6_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmtens.q_2_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpmtens.q_2_LC_6_7_4 .LUT_INIT=16'b1011101110001100;
    LogicCell40 \Lab_UT.didpuu0.didpmtens.q_2_LC_6_7_4  (
            .in0(N__10491),
            .in1(N__13152),
            .in2(N__9795),
            .in3(N__15134),
            .lcout(Lab_UT_di_Mtens_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13500),
            .ce(),
            .sr(N__15880));
    defparam \Lab_UT.dec3.segmentUQ_1_1_LC_6_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dec3.segmentUQ_1_1_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec3.segmentUQ_1_1_LC_6_7_5 .LUT_INIT=16'b0011010111110111;
    LogicCell40 \Lab_UT.dec3.segmentUQ_1_1_LC_6_7_5  (
            .in0(N__15130),
            .in1(N__17005),
            .in2(N__17422),
            .in3(N__15046),
            .lcout(),
            .ltout(Lab_UT_dec3_segmentUQ_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment4_0_bm_LC_6_7_6 .C_ON=1'b0;
    defparam \uu2.un1_segment4_0_bm_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_0_bm_LC_6_7_6 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \uu2.un1_segment4_0_bm_LC_6_7_6  (
            .in0(N__15048),
            .in1(N__17400),
            .in2(N__10380),
            .in3(N__11406),
            .lcout(\uu2.un1_segment4_0_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpmtens.q_RNITG5_1_LC_6_7_7 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmtens.q_RNITG5_1_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpmtens.q_RNITG5_1_LC_6_7_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \Lab_UT.didpuu0.didpmtens.q_RNITG5_1_LC_6_7_7  (
            .in0(N__15132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17004),
            .lcout(N_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIAPHB1_0_5_LC_6_8_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIAPHB1_0_5_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIAPHB1_0_5_LC_6_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIAPHB1_0_5_LC_6_8_0  (
            .in0(N__13771),
            .in1(N__12213),
            .in2(N__12315),
            .in3(N__12838),
            .lcout(\uu2.Z_decfrac105_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNID8KP2_2_LC_6_8_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNID8KP2_2_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNID8KP2_2_LC_6_8_1 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \uu2.w_addr_displaying_RNID8KP2_2_LC_6_8_1  (
            .in0(N__12839),
            .in1(N__11699),
            .in2(N__12156),
            .in3(N__10455),
            .lcout(\uu2.g0_i_o4_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_1_LC_6_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_1_LC_6_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_1_LC_6_8_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_1_LC_6_8_2  (
            .in0(N__17143),
            .in1(N__17080),
            .in2(_gnd_net_),
            .in3(N__10275),
            .lcout(\Lab_UT.didpuu0.ledDisp00.selLedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13495),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dek.det_N_0_a3_LC_6_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dek.det_N_0_a3_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrluu0.dek.det_N_0_a3_LC_6_8_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrluu0.dek.det_N_0_a3_LC_6_8_4  (
            .in0(N__10262),
            .in1(N__10371),
            .in2(N__10320),
            .in3(N__10281),
            .lcout(\Lab_UT.dicSelectLEDdisp ),
            .ltout(\Lab_UT.dicSelectLEDdisp_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_0_LC_6_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_0_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_0_LC_6_8_5 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_0_LC_6_8_5  (
            .in0(N__17079),
            .in1(_gnd_net_),
            .in2(N__10266),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.didpuu0.ledDisp00.selLedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13495),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_2_LC_6_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_2_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_RNO_2_LC_6_8_6 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \Lab_UT.dictrluu0.dicfsm.cState_RNO_2_LC_6_8_6  (
            .in0(N__10263),
            .in1(N__10251),
            .in2(_gnd_net_),
            .in3(N__16569),
            .lcout(),
            .ltout(\Lab_UT.dictrluu0.dicfsm.N_102_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dicfsm.cState_LC_6_8_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_LC_6_8_7 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \Lab_UT.dictrluu0.dicfsm.cState_LC_6_8_7  (
            .in0(N__10245),
            .in1(N__10236),
            .in2(N__10230),
            .in3(N__15921),
            .lcout(Lab_UT_dicRun),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13495),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIAGS21_4_LC_6_9_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIAGS21_4_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIAGS21_4_LC_6_9_0 .LUT_INIT=16'b1010010110101110;
    LogicCell40 \uu2.w_addr_displaying_RNIAGS21_4_LC_6_9_0  (
            .in0(N__13775),
            .in1(N__14462),
            .in2(N__14766),
            .in3(N__13996),
            .lcout(\uu2.un1_segment3_m4_s_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIU2OL2_5_LC_6_9_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIU2OL2_5_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIU2OL2_5_LC_6_9_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIU2OL2_5_LC_6_9_1  (
            .in0(N__13014),
            .in1(N__14510),
            .in2(N__11451),
            .in3(N__10454),
            .lcout(),
            .ltout(\uu2.N_49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI9HV1J_5_LC_6_9_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI9HV1J_5_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI9HV1J_5_LC_6_9_2 .LUT_INIT=16'b0101010001010111;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI9HV1J_5_LC_6_9_2  (
            .in0(N__14472),
            .in1(N__12597),
            .in2(N__10443),
            .in3(N__10395),
            .lcout(\uu2.un1_segment3_m4_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIAH4P4_4_LC_6_9_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIAH4P4_4_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIAH4P4_4_LC_6_9_3 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \uu2.w_addr_displaying_RNIAH4P4_4_LC_6_9_3  (
            .in0(N__10440),
            .in1(N__11619),
            .in2(_gnd_net_),
            .in3(N__11466),
            .lcout(),
            .ltout(\uu2.g0_i_o4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNINK1T81_2_LC_6_9_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNINK1T81_2_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNINK1T81_2_LC_6_9_4 .LUT_INIT=16'b0011011100110010;
    LogicCell40 \uu2.w_addr_displaying_RNINK1T81_2_LC_6_9_4  (
            .in0(N__10434),
            .in1(N__10428),
            .in2(N__10422),
            .in3(N__11478),
            .lcout(\uu2.un1_segment3_m4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep1_RNIMMRIA_LC_6_9_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep1_RNIMMRIA_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_4_rep1_RNIMMRIA_LC_6_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.w_addr_displaying_4_rep1_RNIMMRIA_LC_6_9_5  (
            .in0(N__12666),
            .in1(N__10464),
            .in2(_gnd_net_),
            .in3(N__11364),
            .lcout(\uu2.w_addr_displaying_4_rep1_RNIMMRIAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_6_10_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_6_10_0 .LUT_INIT=16'b1011111110111010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_53_LC_6_10_0  (
            .in0(N__12631),
            .in1(N__14398),
            .in2(N__11607),
            .in3(N__12731),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_53_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_6_10_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_6_10_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_40_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__10515),
            .in2(N__10389),
            .in3(N__11508),
            .lcout(\uu2.mem0.un1_segment3_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_6_rep1_RNI9Q3H_LC_6_10_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_rep1_RNI9Q3H_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_6_rep1_RNI9Q3H_LC_6_10_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uu2.w_addr_displaying_6_rep1_RNI9Q3H_LC_6_10_2  (
            .in0(N__14827),
            .in1(N__15457),
            .in2(_gnd_net_),
            .in3(N__16422),
            .lcout(\uu2.un1_segment4_sn_N_58_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_6_10_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_6_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_52_LC_6_10_3  (
            .in0(N__15747),
            .in1(N__14427),
            .in2(_gnd_net_),
            .in3(N__10527),
            .lcout(\uu2.mem0.un1_segment3_m2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_6_10_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_6_10_4 .LUT_INIT=16'b1011111110111010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_42_LC_6_10_4  (
            .in0(N__12630),
            .in1(N__14397),
            .in2(N__11606),
            .in3(N__12730),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_6_10_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_6_10_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_30_LC_6_10_5  (
            .in0(N__10509),
            .in1(_gnd_net_),
            .in2(N__10503),
            .in3(N__11544),
            .lcout(\uu2.mem0.un1_segment3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec0.un137_segmentUQ_LC_6_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dec0.un137_segmentUQ_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec0.un137_segmentUQ_LC_6_10_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dec0.un137_segmentUQ_LC_6_10_6  (
            .in0(N__14750),
            .in1(N__17246),
            .in2(N__14671),
            .in3(N__15729),
            .lcout(Lab_UT_dec0_un137_segmentUQ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment4_5_am_1_LC_6_10_7 .C_ON=1'b0;
    defparam \uu2.un1_segment4_5_am_1_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_5_am_1_LC_6_10_7 .LUT_INIT=16'b0000001100101010;
    LogicCell40 \uu2.un1_segment4_5_am_1_LC_6_10_7  (
            .in0(N__15730),
            .in1(N__14651),
            .in2(N__17255),
            .in3(N__14751),
            .lcout(\uu2.un1_segment4_5_amZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpmtens.q_RNO_0_2_LC_6_11_0 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmtens.q_RNO_0_2_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpmtens.q_RNO_0_2_LC_6_11_0 .LUT_INIT=16'b0100110001000100;
    LogicCell40 \Lab_UT.didpuu0.didpmtens.q_RNO_0_2_LC_6_11_0  (
            .in0(N__17448),
            .in1(N__15167),
            .in2(N__17063),
            .in3(N__15073),
            .lcout(\Lab_UT.didpuu0.didpmtens.q_5_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment4_1_bm_LC_6_11_1 .C_ON=1'b0;
    defparam \uu2.un1_segment4_1_bm_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_1_bm_LC_6_11_1 .LUT_INIT=16'b0110011010111101;
    LogicCell40 \uu2.un1_segment4_1_bm_LC_6_11_1  (
            .in0(N__15166),
            .in1(N__17054),
            .in2(N__15088),
            .in3(N__17447),
            .lcout(),
            .ltout(\uu2.un1_segment4_1_bmZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIPN54_8_LC_6_11_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIPN54_8_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIPN54_8_LC_6_11_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIPN54_8_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(N__10479),
            .in2(N__10470),
            .in3(N__15248),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_fast_RNIPN54Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI9TKJ4_2_LC_6_11_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI9TKJ4_2_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI9TKJ4_2_LC_6_11_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI9TKJ4_2_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(N__13972),
            .in2(N__10467),
            .in3(N__10581),
            .lcout(\uu2.N_292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIV5694_2_LC_6_11_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIV5694_2_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIV5694_2_LC_6_11_4 .LUT_INIT=16'b1111000000010001;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIV5694_2_LC_6_11_4  (
            .in0(N__10590),
            .in1(N__12868),
            .in2(N__10626),
            .in3(N__12954),
            .lcout(\uu2.w_addr_displaying_fast_RNIV5694Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIHV86_5_LC_6_11_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIHV86_5_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIHV86_5_LC_6_11_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIHV86_5_LC_6_11_5  (
            .in0(N__14568),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14511),
            .lcout(\uu2.N_290_0_i_0 ),
            .ltout(\uu2.N_290_0_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI1BU61_7_LC_6_11_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI1BU61_7_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI1BU61_7_LC_6_11_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI1BU61_7_LC_6_11_6  (
            .in0(N__12795),
            .in1(N__13762),
            .in2(N__10575),
            .in3(N__16278),
            .lcout(),
            .ltout(\uu2.un1_w_addr_displaying_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI90195_7_LC_6_11_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI90195_7_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI90195_7_LC_6_11_7 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \uu2.w_addr_displaying_RNI90195_7_LC_6_11_7  (
            .in0(N__16279),
            .in1(N__10572),
            .in2(N__10566),
            .in3(N__16482),
            .lcout(\uu2.un1_w_addr_displaying_inv_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_6_12_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_6_12_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_51_LC_6_12_1  (
            .in0(N__13770),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12812),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_6_12_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_6_12_2 .LUT_INIT=16'b1000000011111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_39_LC_6_12_2  (
            .in0(N__12224),
            .in1(N__12291),
            .in2(N__10563),
            .in3(N__11595),
            .lcout(\uu2.mem0.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIAPHB1_5_LC_6_12_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIAPHB1_5_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIAPHB1_5_LC_6_12_3 .LUT_INIT=16'b1011111101111111;
    LogicCell40 \uu2.w_addr_displaying_RNIAPHB1_5_LC_6_12_3  (
            .in0(N__13769),
            .in1(N__12223),
            .in2(N__12305),
            .in3(N__12811),
            .lcout(\uu2.un1_segment3_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_5_LC_6_12_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_LC_6_12_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_LC_6_12_5 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \uu2.w_addr_displaying_5_LC_6_12_5  (
            .in0(N__12292),
            .in1(_gnd_net_),
            .in2(N__13916),
            .in3(N__16103),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_5C_net ),
            .ce(),
            .sr(N__15854));
    defparam \uu2.w_addr_displaying_3_LC_6_12_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_LC_6_12_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.w_addr_displaying_3_LC_6_12_6  (
            .in0(N__12813),
            .in1(N__15492),
            .in2(_gnd_net_),
            .in3(N__16102),
            .lcout(\uu2.w_addr_displayingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_5C_net ),
            .ce(),
            .sr(N__15854));
    defparam \uu2.w_addr_displaying_0_rep1_RNIUUGB1_LC_6_12_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_RNIUUGB1_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_0_rep1_RNIUUGB1_LC_6_12_7 .LUT_INIT=16'b0001000000000100;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_RNIUUGB1_LC_6_12_7  (
            .in0(N__11460),
            .in1(N__12810),
            .in2(N__13780),
            .in3(N__14312),
            .lcout(\uu2.un1_segment4_sn_N_38_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment4_2_bm_LC_6_13_0 .C_ON=1'b0;
    defparam \uu2.un1_segment4_2_bm_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_2_bm_LC_6_13_0 .LUT_INIT=16'b0011110101010111;
    LogicCell40 \uu2.un1_segment4_2_bm_LC_6_13_0  (
            .in0(N__14744),
            .in1(N__17248),
            .in2(N__14674),
            .in3(N__15732),
            .lcout(\uu2.un1_segment4_2_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.g1_LC_6_13_1 .C_ON=1'b0;
    defparam \uu2.g1_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \uu2.g1_LC_6_13_1 .LUT_INIT=16'b1111101101111100;
    LogicCell40 \uu2.g1_LC_6_13_1  (
            .in0(N__15733),
            .in1(N__14745),
            .in2(N__17256),
            .in3(N__14664),
            .lcout(\uu2.gZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment4_5_bm_LC_6_13_2 .C_ON=1'b0;
    defparam \uu2.un1_segment4_5_bm_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_5_bm_LC_6_13_2 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \uu2.un1_segment4_5_bm_LC_6_13_2  (
            .in0(N__14743),
            .in1(N__17247),
            .in2(N__14673),
            .in3(N__15731),
            .lcout(\uu2.un1_segment4_5_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_3_LC_6_13_3 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_3_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_3_LC_6_13_3 .LUT_INIT=16'b0111011111011101;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_RNO_0_3_LC_6_13_3  (
            .in0(N__15734),
            .in1(N__14747),
            .in2(_gnd_net_),
            .in3(N__17253),
            .lcout(\Lab_UT.didpuu0.didpsones.N_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_RNI0GG11_3_LC_6_13_4 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_RNI0GG11_3_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpsones.q_RNI0GG11_3_LC_6_13_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_RNI0GG11_3_LC_6_13_4  (
            .in0(N__14746),
            .in1(_gnd_net_),
            .in2(N__14675),
            .in3(N__17252),
            .lcout(\Lab_UT.didpuu0.didpsones.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMU_0_LC_6_13_5 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMU_0_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMU_0_LC_6_13_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMU_0_LC_6_13_5  (
            .in0(N__17093),
            .in1(N__14191),
            .in2(_gnd_net_),
            .in3(N__14748),
            .lcout(),
            .ltout(\Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMUZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIEH0Q1_1_LC_6_13_6 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIEH0Q1_1_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIEH0Q1_1_LC_6_13_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNIEH0Q1_1_LC_6_13_6  (
            .in0(N__17150),
            .in1(_gnd_net_),
            .in2(N__10614),
            .in3(N__10596),
            .lcout(led_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJ_0_LC_6_13_7 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJ_0_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJ_0_LC_6_13_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJ_0_LC_6_13_7  (
            .in0(N__17094),
            .in1(N__16970),
            .in2(_gnd_net_),
            .in3(N__15188),
            .lcout(\Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_LC_7_2_0 .C_ON=1'b1;
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_LC_7_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.un1_bitcount_cry_0_c_LC_7_2_0  (
            .in0(_gnd_net_),
            .in1(N__10632),
            .in2(N__10701),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_2_0_),
            .carryout(\buart.Z_tx.un1_bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_1_LC_7_2_1 .C_ON=1'b1;
    defparam \buart.Z_tx.bitcount_1_LC_7_2_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_1_LC_7_2_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_7_2_1  (
            .in0(N__11164),
            .in1(N__10755),
            .in2(N__10731),
            .in3(N__10776),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(\buart.Z_tx.un1_bitcount_cry_0 ),
            .carryout(\buart.Z_tx.un1_bitcount_cry_1 ),
            .clk(N__13543),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_2_LC_7_2_2 .C_ON=1'b1;
    defparam \buart.Z_tx.bitcount_2_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_2_LC_7_2_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_7_2_2  (
            .in0(N__11165),
            .in1(N__10761),
            .in2(N__10749),
            .in3(N__10773),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.un1_bitcount_cry_1 ),
            .carryout(\buart.Z_tx.un1_bitcount_cry_2 ),
            .clk(N__13543),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_3_LC_7_2_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_7_2_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_3_LC_7_2_3 .LUT_INIT=16'b1101110111101110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_7_2_3  (
            .in0(N__10770),
            .in1(N__11166),
            .in2(_gnd_net_),
            .in3(N__10764),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13543),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIM5O32_2_LC_7_2_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIM5O32_2_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIM5O32_2_LC_7_2_4 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \buart.Z_tx.bitcount_RNIM5O32_2_LC_7_2_4  (
            .in0(N__10668),
            .in1(_gnd_net_),
            .in2(N__10813),
            .in3(N__10748),
            .lcout(\buart.Z_tx.bitcount_RNIM5O32Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIL4O32_1_LC_7_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIL4O32_1_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIL4O32_1_LC_7_2_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIL4O32_1_LC_7_2_5  (
            .in0(N__10730),
            .in1(N__10801),
            .in2(_gnd_net_),
            .in3(N__10667),
            .lcout(\buart.Z_tx.bitcount_RNIL4O32Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_7_2_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_7_2_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_tx.bitcount_RNIQOQA1_3_LC_7_2_6  (
            .in0(N__10744),
            .in1(N__10726),
            .in2(N__10716),
            .in3(N__10695),
            .lcout(buart__tx_uart_busy_0),
            .ltout(buart__tx_uart_busy_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_RNO_LC_7_2_7 .C_ON=1'b0;
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_RNO_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_RNO_LC_7_2_7 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \buart.Z_tx.un1_bitcount_cry_0_c_RNO_LC_7_2_7  (
            .in0(N__10696),
            .in1(_gnd_net_),
            .in2(N__10677),
            .in3(N__10666),
            .lcout(\buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_8_LC_7_3_7 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_7_3_7 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_8_LC_7_3_7 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.l_count_8_LC_7_3_7  (
            .in0(N__12101),
            .in1(N__12009),
            .in2(_gnd_net_),
            .in3(N__12077),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13537),
            .ce(),
            .sr(N__15890));
    defparam \resetGen.reset_count_RNITEEC1_2_LC_7_4_0 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNITEEC1_2_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNITEEC1_2_LC_7_4_0 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \resetGen.reset_count_RNITEEC1_2_LC_7_4_0  (
            .in0(N__10905),
            .in1(N__10891),
            .in2(_gnd_net_),
            .in3(N__10823),
            .lcout(\resetGen.N_117 ),
            .ltout(\resetGen.N_117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_7_4_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_7_4_1 .LUT_INIT=16'b0000000011001110;
    LogicCell40 \resetGen.reset_count_4_LC_7_4_1  (
            .in0(N__10955),
            .in1(N__10880),
            .in2(N__10941),
            .in3(N__10851),
            .lcout(\resetGen.reset_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13530),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_7_4_2 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_7_4_2 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \resetGen.reset_count_1_LC_7_4_2  (
            .in0(N__10849),
            .in1(N__10878),
            .in2(N__10911),
            .in3(N__10893),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13530),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_7_4_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_7_4_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_7_4_3 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \resetGen.reset_count_0_LC_7_4_3  (
            .in0(N__10877),
            .in1(N__10907),
            .in2(_gnd_net_),
            .in3(N__10848),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13530),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_7_4_4 .C_ON=1'b0;
    defparam \resetGen.rst_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_7_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_7_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10876),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13530),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNO_0_2_LC_7_4_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_2_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_2_LC_7_4_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \resetGen.reset_count_RNO_0_2_LC_7_4_6  (
            .in0(N__10906),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10892),
            .lcout(),
            .ltout(\resetGen.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_7_4_7 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_7_4_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_7_4_7 .LUT_INIT=16'b0000000010101001;
    LogicCell40 \resetGen.reset_count_2_LC_7_4_7  (
            .in0(N__10824),
            .in1(N__10879),
            .in2(N__10854),
            .in3(N__10850),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13530),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_10__un382_ci_8_1_LC_7_5_0 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_10__un382_ci_8_1_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_10__un382_ci_8_1_LC_7_5_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_10__un382_ci_8_1_LC_7_5_0  (
            .in0(N__12131),
            .in1(N__11952),
            .in2(N__12054),
            .in3(N__11977),
            .lcout(\uu2.vbuf_count.un382_ci_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_7__un349_ci_0_LC_7_5_1 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_7__un349_ci_0_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_7__un349_ci_0_LC_7_5_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_7__un349_ci_0_LC_7_5_1  (
            .in0(N__11978),
            .in1(N__12052),
            .in2(_gnd_net_),
            .in3(N__11953),
            .lcout(\uu2.un349_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIQF5F5_4_LC_7_5_2 .C_ON=1'b0;
    defparam \uu2.l_count_RNIQF5F5_4_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIQF5F5_4_LC_7_5_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.l_count_RNIQF5F5_4_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(N__10814),
            .in2(_gnd_net_),
            .in3(N__11913),
            .lcout(vbuf_tx_data_rdy),
            .ltout(vbuf_tx_data_rdy_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIU80H5_4_LC_7_5_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNIU80H5_4_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIU80H5_4_LC_7_5_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uu2.l_count_RNIU80H5_4_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11355),
            .in3(N__15920),
            .lcout(\uu2.vbuf_tx_data_rdy_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_4_LC_7_5_4 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_4_LC_7_5_4 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \uu2.l_count_4_LC_7_5_4  (
            .in0(N__12053),
            .in1(N__12017),
            .in2(_gnd_net_),
            .in3(N__11914),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13525),
            .ce(),
            .sr(N__15886));
    defparam \uu2.r_addr_1_LC_7_5_6 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_7_5_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.r_addr_1_LC_7_5_6  (
            .in0(N__11279),
            .in1(N__11304),
            .in2(_gnd_net_),
            .in3(N__11162),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13525),
            .ce(),
            .sr(N__15886));
    defparam \uu2.r_addr_2_LC_7_6_2 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_7_6_2 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_2_LC_7_6_2  (
            .in0(N__11305),
            .in1(N__11272),
            .in2(N__11103),
            .in3(N__11163),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13518),
            .ce(),
            .sr(N__15884));
    defparam \Lab_UT.didpuu0.didpmtens.q_0_LC_7_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmtens.q_0_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpmtens.q_0_LC_7_7_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \Lab_UT.didpuu0.didpmtens.q_0_LC_7_7_2  (
            .in0(N__13215),
            .in1(N__13183),
            .in2(_gnd_net_),
            .in3(N__17420),
            .lcout(Lab_UT_di_Mtens_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13511),
            .ce(),
            .sr(N__15883));
    defparam \uu2.un1_segment4_2_am_LC_7_7_4 .C_ON=1'b0;
    defparam \uu2.un1_segment4_2_am_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_2_am_LC_7_7_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uu2.un1_segment4_2_am_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__12240),
            .in2(_gnd_net_),
            .in3(N__12872),
            .lcout(\uu2.un1_segment4_2_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.sec_clk_LC_7_7_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.sec_clk_LC_7_7_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.sec_clk_LC_7_7_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.secuu0.sec_clk_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__11076),
            .in2(_gnd_net_),
            .in3(N__16537),
            .lcout(Lab_UT_l_oneSecPluse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13511),
            .ce(),
            .sr(N__15883));
    defparam \Lab_UT.secuu0.delay_line_1_LC_7_7_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.delay_line_1_LC_7_7_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.delay_line_1_LC_7_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.secuu0.delay_line_1_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10995),
            .lcout(\Lab_UT.secuu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13511),
            .ce(),
            .sr(N__15883));
    defparam \Lab_UT.didpuu0.didpmtens.q_1_LC_7_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmtens.q_1_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpmtens.q_1_LC_7_8_0 .LUT_INIT=16'b0100011001001100;
    LogicCell40 \Lab_UT.didpuu0.didpmtens.q_1_LC_7_8_0  (
            .in0(N__13151),
            .in1(N__17045),
            .in2(N__11418),
            .in3(N__17419),
            .lcout(Lab_UT_di_Mtens_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13502),
            .ce(),
            .sr(N__15879));
    defparam \Lab_UT.didpuu0.didpmtens.q_RNO_0_1_LC_7_8_1 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmtens.q_RNO_0_1_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpmtens.q_RNO_0_1_LC_7_8_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.didpuu0.didpmtens.q_RNO_0_1_LC_7_8_1  (
            .in0(N__17417),
            .in1(N__15051),
            .in2(_gnd_net_),
            .in3(N__15137),
            .lcout(\Lab_UT.didpuu0.didpmtens.N_122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec3.segmentUQ_0_o2_5_LC_7_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dec3.segmentUQ_0_o2_5_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec3.segmentUQ_0_o2_5_LC_7_8_2 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \Lab_UT.dec3.segmentUQ_0_o2_5_LC_7_8_2  (
            .in0(N__15135),
            .in1(N__17043),
            .in2(_gnd_net_),
            .in3(N__17415),
            .lcout(),
            .ltout(N_84_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment4_0_am_LC_7_8_3 .C_ON=1'b0;
    defparam \uu2.un1_segment4_0_am_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_0_am_LC_7_8_3 .LUT_INIT=16'b1101110001110011;
    LogicCell40 \uu2.un1_segment4_0_am_LC_7_8_3  (
            .in0(N__17416),
            .in1(N__15050),
            .in2(N__11409),
            .in3(N__11405),
            .lcout(),
            .ltout(\uu2.un1_segment4_0_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIK7I7_2_LC_7_8_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIK7I7_2_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIK7I7_2_LC_7_8_4 .LUT_INIT=16'b0011001101000111;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIK7I7_2_LC_7_8_4  (
            .in0(N__11394),
            .in1(N__12962),
            .in2(N__11388),
            .in3(N__12988),
            .lcout(),
            .ltout(\uu2.un1_segment4_8_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep1_RNI6JSF4_LC_7_8_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep1_RNI6JSF4_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_4_rep1_RNI6JSF4_LC_7_8_5 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \uu2.w_addr_displaying_4_rep1_RNI6JSF4_LC_7_8_5  (
            .in0(N__11385),
            .in1(N__14822),
            .in2(N__11373),
            .in3(N__11370),
            .lcout(\uu2.N_286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec3.un75_segmentUQ_i_i_o2_LC_7_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dec3.un75_segmentUQ_i_i_o2_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec3.un75_segmentUQ_i_i_o2_LC_7_8_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.dec3.un75_segmentUQ_i_i_o2_LC_7_8_6  (
            .in0(N__15136),
            .in1(N__17044),
            .in2(_gnd_net_),
            .in3(N__17418),
            .lcout(),
            .ltout(\Lab_UT.N_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpmtens.q_3_LC_7_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmtens.q_3_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpmtens.q_3_LC_7_8_7 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \Lab_UT.didpuu0.didpmtens.q_3_LC_7_8_7  (
            .in0(N__13184),
            .in1(N__13214),
            .in2(N__11358),
            .in3(N__15052),
            .lcout(Lab_UT_di_Mtens_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13502),
            .ce(),
            .sr(N__15879));
    defparam \uu2.w_addr_displaying_fast_RNIK9D9_2_LC_7_9_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIK9D9_2_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIK9D9_2_LC_7_9_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIK9D9_2_LC_7_9_0  (
            .in0(N__12952),
            .in1(N__14554),
            .in2(_gnd_net_),
            .in3(N__13060),
            .lcout(\uu2.un1_segment4_sn_N_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNILAD9_2_LC_7_9_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNILAD9_2_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNILAD9_2_LC_7_9_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNILAD9_2_LC_7_9_1  (
            .in0(N__14555),
            .in1(N__12953),
            .in2(_gnd_net_),
            .in3(N__12989),
            .lcout(),
            .ltout(\uu2.g0_i_o4_0_a8_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_5_rep1_RNIVO2E1_LC_7_9_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_rep1_RNIVO2E1_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_5_rep1_RNIVO2E1_LC_7_9_2 .LUT_INIT=16'b0101010100010101;
    LogicCell40 \uu2.w_addr_displaying_5_rep1_RNIVO2E1_LC_7_9_2  (
            .in0(N__12924),
            .in1(N__13851),
            .in2(N__11469),
            .in3(N__16473),
            .lcout(\uu2.w_addr_displaying_5_rep1_RNIVO2EZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_4_LC_7_9_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_4_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_4_LC_7_9_3 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.w_addr_displaying_fast_4_LC_7_9_3  (
            .in0(N__15292),
            .in1(_gnd_net_),
            .in2(N__16092),
            .in3(N__12990),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_4C_net ),
            .ce(),
            .sr(N__15850));
    defparam \uu2.w_addr_displaying_fast_6_LC_7_9_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_6_LC_7_9_4 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_fast_6_LC_7_9_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uu2.w_addr_displaying_fast_6_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__16049),
            .in2(N__12585),
            .in3(N__14556),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_4C_net ),
            .ce(),
            .sr(N__15850));
    defparam \uu2.w_addr_displaying_8_rep1_LC_7_9_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_rep1_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_rep1_LC_7_9_5 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_8_rep1_LC_7_9_5  (
            .in0(N__13852),
            .in1(N__16059),
            .in2(N__15306),
            .in3(N__15369),
            .lcout(\uu2.w_addr_displaying_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_4C_net ),
            .ce(),
            .sr(N__15850));
    defparam \uu2.w_addr_displaying_8_rep1_RNIN6OC_LC_7_9_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_rep1_RNIN6OC_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_8_rep1_RNIN6OC_LC_7_9_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uu2.w_addr_displaying_8_rep1_RNIN6OC_LC_7_9_6  (
            .in0(N__13826),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14887),
            .lcout(\uu2.N_315_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_7_rep1_LC_7_9_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_rep1_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_rep1_LC_7_9_7 .LUT_INIT=16'b1010101001101010;
    LogicCell40 \uu2.w_addr_displaying_7_rep1_LC_7_9_7  (
            .in0(N__14888),
            .in1(N__16058),
            .in2(N__13913),
            .in3(N__14013),
            .lcout(\uu2.w_addr_displaying_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_4C_net ),
            .ce(),
            .sr(N__15850));
    defparam \uu2.w_addr_displaying_2_rep1_RNIQ3R01_LC_7_10_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_RNIQ3R01_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_2_rep1_RNIQ3R01_LC_7_10_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_RNIQ3R01_LC_7_10_0  (
            .in0(N__15458),
            .in1(N__14307),
            .in2(N__15552),
            .in3(N__16365),
            .lcout(\uu2.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep2_RNI5R4M_LC_7_10_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep2_RNI5R4M_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_4_rep2_RNI5R4M_LC_7_10_1 .LUT_INIT=16'b0100010010011001;
    LogicCell40 \uu2.w_addr_displaying_4_rep2_RNI5R4M_LC_7_10_1  (
            .in0(N__14308),
            .in1(N__11685),
            .in2(_gnd_net_),
            .in3(N__15551),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_1_1_3_tz_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIDUPM1_2_LC_7_10_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIDUPM1_2_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIDUPM1_2_LC_7_10_2 .LUT_INIT=16'b1110111110011111;
    LogicCell40 \uu2.w_addr_displaying_RNIDUPM1_2_LC_7_10_2  (
            .in0(N__11686),
            .in1(N__12834),
            .in2(N__11442),
            .in3(N__14999),
            .lcout(\uu2.bitmap_pmux_1_1_3_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI50L01_2_LC_7_10_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI50L01_2_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI50L01_2_LC_7_10_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI50L01_2_LC_7_10_4  (
            .in0(N__11687),
            .in1(N__16184),
            .in2(_gnd_net_),
            .in3(N__15000),
            .lcout(\uu2.N_111 ),
            .ltout(\uu2.N_111_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_5__un436_ci_0_a2_LC_7_10_5 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_5__un436_ci_0_a2_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_5__un436_ci_0_a2_LC_7_10_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uu2.vbuf_w_addr_displaying.counter_gen_label_5__un436_ci_0_a2_LC_7_10_5  (
            .in0(N__12835),
            .in1(_gnd_net_),
            .in2(N__11523),
            .in3(N__13757),
            .lcout(\uu2.un436_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_LC_7_10_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_LC_7_10_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.w_addr_displaying_4_LC_7_10_6  (
            .in0(N__13758),
            .in1(N__15291),
            .in2(_gnd_net_),
            .in3(N__16083),
            .lcout(\uu2.w_addr_displayingZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__15852));
    defparam \uu2.w_addr_displaying_fast_2_LC_7_10_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_2_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_2_LC_7_10_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_fast_2_LC_7_10_7  (
            .in0(N__16082),
            .in1(N__15001),
            .in2(N__16199),
            .in3(N__12961),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__15852));
    defparam \uu2.w_addr_displaying_5_rep1_RNI50LS_LC_7_11_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_rep1_RNI50LS_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_5_rep1_RNI50LS_LC_7_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_5_rep1_RNI50LS_LC_7_11_0  (
            .in0(N__16421),
            .in1(N__15459),
            .in2(N__14902),
            .in3(N__16472),
            .lcout(),
            .ltout(\uu2.un1_segment4_sn_N_36_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_5_rep1_RNIMG8P2_LC_7_11_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_rep1_RNIMG8P2_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_5_rep1_RNIMG8P2_LC_7_11_1 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \uu2.w_addr_displaying_5_rep1_RNIMG8P2_LC_7_11_1  (
            .in0(N__16547),
            .in1(N__16570),
            .in2(N__11520),
            .in3(N__11517),
            .lcout(\uu2.N_2150_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_7_11_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_7_11_2 .LUT_INIT=16'b0001001100010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_54_LC_7_11_2  (
            .in0(N__14386),
            .in1(N__12618),
            .in2(N__11599),
            .in3(N__12715),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIKR5D1_6_LC_7_11_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIKR5D1_6_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIKR5D1_6_LC_7_11_3 .LUT_INIT=16'b0001001111111111;
    LogicCell40 \uu2.w_addr_displaying_RNIKR5D1_6_LC_7_11_3  (
            .in0(N__12222),
            .in1(N__11502),
            .in2(N__12575),
            .in3(N__13983),
            .lcout(),
            .ltout(\uu2.g2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_rep1_RNIN998E_LC_7_11_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_RNIN998E_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_0_rep1_RNIN998E_LC_7_11_4 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_RNIN998E_LC_7_11_4  (
            .in0(N__11496),
            .in1(N__11490),
            .in2(N__11481),
            .in3(N__13089),
            .lcout(\uu2.N_299_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_7_11_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_7_11_5 .LUT_INIT=16'b0001000101010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_43_LC_7_11_5  (
            .in0(N__12617),
            .in1(N__14385),
            .in2(N__12729),
            .in3(N__11586),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIUCHB1_3_LC_7_11_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIUCHB1_3_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIUCHB1_3_LC_7_11_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIUCHB1_3_LC_7_11_6  (
            .in0(N__15480),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12837),
            .lcout(\uu2.un15_w_data_displaying_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec2.segmentUQ_2_LC_7_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dec2.segmentUQ_2_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec2.segmentUQ_2_LC_7_12_0 .LUT_INIT=16'b0010111111111011;
    LogicCell40 \Lab_UT.dec2.segmentUQ_2_LC_7_12_0  (
            .in0(N__16670),
            .in1(N__16859),
            .in2(N__16965),
            .in3(N__16721),
            .lcout(L3_segment3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpmones.q_esr_3_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmones.q_esr_3_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpmones.q_esr_3_LC_7_12_1 .LUT_INIT=16'b0110100011110000;
    LogicCell40 \Lab_UT.didpuu0.didpmones.q_esr_3_LC_7_12_1  (
            .in0(N__16863),
            .in1(N__16953),
            .in2(N__16743),
            .in3(N__16674),
            .lcout(Lab_UT_di_Mones_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13488),
            .ce(N__11865),
            .sr(N__15887));
    defparam \uu2.segment3_m_1_6_LC_7_12_2 .C_ON=1'b0;
    defparam \uu2.segment3_m_1_6_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \uu2.segment3_m_1_6_LC_7_12_2 .LUT_INIT=16'b1110111101111100;
    LogicCell40 \uu2.segment3_m_1_6_LC_7_12_2  (
            .in0(N__16672),
            .in1(N__16861),
            .in2(N__16964),
            .in3(N__16720),
            .lcout(),
            .ltout(\uu2.segment3_m_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_7_rep1_RNIA86H1_LC_7_12_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_rep1_RNIA86H1_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_7_rep1_RNIA86H1_LC_7_12_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.w_addr_displaying_7_rep1_RNIA86H1_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11538),
            .in3(N__14892),
            .lcout(),
            .ltout(\uu2.segment3_m_2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIE28D2_4_LC_7_12_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIE28D2_4_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIE28D2_4_LC_7_12_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \uu2.w_addr_displaying_RNIE28D2_4_LC_7_12_4  (
            .in0(N__13763),
            .in1(N__12794),
            .in2(N__11535),
            .in3(N__13973),
            .lcout(\uu2.segment3_m_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment4_4_bm_LC_7_12_5 .C_ON=1'b0;
    defparam \uu2.un1_segment4_4_bm_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_4_bm_LC_7_12_5 .LUT_INIT=16'b1110000011111011;
    LogicCell40 \uu2.un1_segment4_4_bm_LC_7_12_5  (
            .in0(N__16860),
            .in1(N__16946),
            .in2(N__16742),
            .in3(N__16671),
            .lcout(\uu2.un1_segment4_4_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment4_4_am_LC_7_12_6 .C_ON=1'b0;
    defparam \uu2.un1_segment4_4_am_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_4_am_LC_7_12_6 .LUT_INIT=16'b1101111101110001;
    LogicCell40 \uu2.un1_segment4_4_am_LC_7_12_6  (
            .in0(N__16673),
            .in1(N__16862),
            .in2(N__16963),
            .in3(N__16716),
            .lcout(),
            .ltout(\uu2.un1_segment4_4_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNICB763_0_LC_7_12_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNICB763_0_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNICB763_0_LC_7_12_7 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \uu2.w_addr_displaying_fast_RNICB763_0_LC_7_12_7  (
            .in0(N__15249),
            .in1(N__11532),
            .in2(N__11526),
            .in3(N__15944),
            .lcout(\uu2.un1_segment4_9_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_7_13_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_7_13_0 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_23_LC_7_13_0  (
            .in0(N__12571),
            .in1(N__11736),
            .in2(N__12483),
            .in3(N__16285),
            .lcout(\uu2.mem0.G_14_0_a6_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_7_13_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_7_13_1 .LUT_INIT=16'b1101101111110111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_36_LC_7_13_1  (
            .in0(N__12799),
            .in1(N__11662),
            .in2(N__11730),
            .in3(N__14993),
            .lcout(\uu2.mem0.bitmap_pmux_1_1_2_tz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI83L01_2_LC_7_13_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI83L01_2_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI83L01_2_LC_7_13_2 .LUT_INIT=16'b0101010111111010;
    LogicCell40 \uu2.w_addr_displaying_RNI83L01_2_LC_7_13_2  (
            .in0(N__13765),
            .in1(_gnd_net_),
            .in2(N__11684),
            .in3(N__16175),
            .lcout(\uu2.bitmap_pmux_1_1_2_tz_1_0 ),
            .ltout(\uu2.bitmap_pmux_1_1_2_tz_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_7_13_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_7_13_3 .LUT_INIT=16'b1101101111110111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_45_LC_7_13_3  (
            .in0(N__12798),
            .in1(N__11661),
            .in2(N__11721),
            .in3(N__14992),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_1_1_2_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_7_13_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_7_13_4 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_33_LC_7_13_4  (
            .in0(N__12570),
            .in1(_gnd_net_),
            .in2(N__11718),
            .in3(N__16284),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_LC_7_13_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_7_13_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_displaying_2_LC_7_13_5  (
            .in0(N__16176),
            .in1(N__11663),
            .in2(N__16104),
            .in3(N__14994),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2C_net ),
            .ce(),
            .sr(N__15857));
    defparam \uu2.w_addr_displaying_RNI8NHB1_2_LC_7_13_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8NHB1_2_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8NHB1_2_LC_7_13_6 .LUT_INIT=16'b0000000010110101;
    LogicCell40 \uu2.w_addr_displaying_RNI8NHB1_2_LC_7_13_6  (
            .in0(N__13764),
            .in1(N__12797),
            .in2(N__11683),
            .in3(N__16283),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_RNI8NHB1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI18582_8_LC_7_13_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI18582_8_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI18582_8_LC_7_13_7 .LUT_INIT=16'b0011001010111010;
    LogicCell40 \uu2.w_addr_displaying_RNI18582_8_LC_7_13_7  (
            .in0(N__13020),
            .in1(N__12569),
            .in2(N__11622),
            .in3(N__13997),
            .lcout(\uu2.w_addr_displaying_RNI18582Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec2.un152_segmentUQ_1_LC_7_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dec2.un152_segmentUQ_1_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec2.un152_segmentUQ_1_LC_7_14_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dec2.un152_segmentUQ_1_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__16754),
            .in2(_gnd_net_),
            .in3(N__16939),
            .lcout(\Lab_UT.un152_segmentUQ_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI89GK1_2_LC_8_3_0 .C_ON=1'b0;
    defparam \uu2.l_count_RNI89GK1_2_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI89GK1_2_LC_8_3_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uu2.l_count_RNI89GK1_2_LC_8_3_0  (
            .in0(N__11955),
            .in1(N__11841),
            .in2(N__12078),
            .in3(N__11821),
            .lcout(\uu2.un3_r_clk_en_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_2_LC_8_3_1 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_2_LC_8_3_1 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uu2.l_count_2_LC_8_3_1  (
            .in0(N__11783),
            .in1(N__11825),
            .in2(N__11849),
            .in3(N__11921),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13544),
            .ce(),
            .sr(N__15893));
    defparam \uu2.l_count_0_LC_8_3_2 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_0_LC_8_3_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uu2.l_count_0_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__11822),
            .in2(_gnd_net_),
            .in3(N__11919),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13544),
            .ce(),
            .sr(N__15893));
    defparam \uu2.l_count_3_LC_8_3_3 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_3_LC_8_3_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.l_count_3_LC_8_3_3  (
            .in0(N__11784),
            .in1(N__11848),
            .in2(N__11802),
            .in3(N__11826),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13544),
            .ce(),
            .sr(N__15893));
    defparam \uu2.vbuf_count.counter_gen_label_4__un316_ci_LC_8_3_4 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un316_ci_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un316_ci_LC_8_3_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un316_ci_LC_8_3_4  (
            .in0(N__11823),
            .in1(N__11798),
            .in2(N__11850),
            .in3(N__11781),
            .lcout(\uu2.un316_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_1_LC_8_3_7 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_8_3_7 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_1_LC_8_3_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.l_count_1_LC_8_3_7  (
            .in0(N__11782),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11824),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13544),
            .ce(),
            .sr(N__15893));
    defparam \uu2.l_count_RNI89GK1_3_LC_8_4_0 .C_ON=1'b0;
    defparam \uu2.l_count_RNI89GK1_3_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI89GK1_3_LC_8_4_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uu2.l_count_RNI89GK1_3_LC_8_4_0  (
            .in0(N__11975),
            .in1(N__11797),
            .in2(N__12132),
            .in3(N__11780),
            .lcout(\uu2.un3_r_clk_en_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI626E_10_LC_8_4_2 .C_ON=1'b0;
    defparam \uu2.l_count_RNI626E_10_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI626E_10_LC_8_4_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uu2.l_count_RNI626E_10_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(N__11879),
            .in2(_gnd_net_),
            .in3(N__12112),
            .lcout(),
            .ltout(\uu2.un3_r_clk_en_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI0NA44_4_LC_8_4_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNI0NA44_4_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI0NA44_4_LC_8_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI0NA44_4_LC_8_4_3  (
            .in0(N__12039),
            .in1(N__11763),
            .in2(N__11757),
            .in3(N__11754),
            .lcout(uu2_un3_r_clk_en_0),
            .ltout(uu2_un3_r_clk_en_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_5_LC_8_4_4 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_5_LC_8_4_4 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \uu2.l_count_5_LC_8_4_4  (
            .in0(N__11976),
            .in1(N__12008),
            .in2(N__12144),
            .in3(N__12040),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13538),
            .ce(),
            .sr(N__15892));
    defparam \uu2.l_count_7_LC_8_4_5 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_7_LC_8_4_5 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu2.l_count_7_LC_8_4_5  (
            .in0(N__12006),
            .in1(N__12130),
            .in2(N__12141),
            .in3(N__11918),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13538),
            .ce(),
            .sr(N__15892));
    defparam \uu2.l_count_9_LC_8_4_6 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_9_LC_8_4_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.l_count_9_LC_8_4_6  (
            .in0(N__12076),
            .in1(N__12007),
            .in2(N__12102),
            .in3(N__12114),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13538),
            .ce(),
            .sr(N__15892));
    defparam \uu2.vbuf_count.counter_gen_label_10__un382_ci_LC_8_4_7 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_10__un382_ci_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_10__un382_ci_LC_8_4_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_10__un382_ci_LC_8_4_7  (
            .in0(N__12113),
            .in1(N__12097),
            .in2(N__12016),
            .in3(N__12075),
            .lcout(\uu2.un382_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_6_LC_8_5_4 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_6_LC_8_5_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.l_count_6_LC_8_5_4  (
            .in0(N__12048),
            .in1(N__11954),
            .in2(N__12021),
            .in3(N__11979),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13531),
            .ce(),
            .sr(N__15889));
    defparam \uu2.l_count_10_LC_8_5_6 .C_ON=1'b0;
    defparam \uu2.l_count_10_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_10_LC_8_5_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \uu2.l_count_10_LC_8_5_6  (
            .in0(N__11928),
            .in1(N__11880),
            .in2(_gnd_net_),
            .in3(N__11920),
            .lcout(\uu2.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13531),
            .ce(),
            .sr(N__15889));
    defparam \Lab_UT.didpuu0.didpstens.q_RNIL3BL3_1_LC_8_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpstens.q_RNIL3BL3_1_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpstens.q_RNIL3BL3_1_LC_8_7_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.didpuu0.didpstens.q_RNIL3BL3_1_LC_8_7_0  (
            .in0(N__13177),
            .in1(N__17325),
            .in2(N__13244),
            .in3(N__15635),
            .lcout(\Lab_UT.didpuu0.countEnMones ),
            .ltout(\Lab_UT.didpuu0.countEnMones_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpmones.q_esr_RNO_0_3_LC_8_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmones.q_esr_RNO_0_3_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpmones.q_esr_RNO_0_3_LC_8_7_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.didpuu0.didpmones.q_esr_RNO_0_3_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11868),
            .in3(N__15918),
            .lcout(\Lab_UT.didpuu0.didpmones.countEnMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpstens.q_1_LC_8_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpstens.q_1_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpstens.q_1_LC_8_7_2 .LUT_INIT=16'b0100011011001100;
    LogicCell40 \Lab_UT.didpuu0.didpstens.q_1_LC_8_7_2  (
            .in0(N__13179),
            .in1(N__17326),
            .in2(N__13245),
            .in3(N__15637),
            .lcout(Lab_UT_di_Stens_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13519),
            .ce(),
            .sr(N__15885));
    defparam \Lab_UT.didpuu0.didpstens.q_0_LC_8_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpstens.q_0_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpstens.q_0_LC_8_7_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.didpuu0.didpstens.q_0_LC_8_7_3  (
            .in0(N__15636),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13178),
            .lcout(Lab_UT_di_Stens_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13519),
            .ce(),
            .sr(N__15885));
    defparam \Lab_UT.didpuu0.didpsones.q_RNIHCAV1_0_LC_8_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_RNIHCAV1_0_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpsones.q_RNIHCAV1_0_LC_8_7_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_RNIHCAV1_0_LC_8_7_4  (
            .in0(N__15690),
            .in1(N__12917),
            .in2(_gnd_net_),
            .in3(N__13306),
            .lcout(\Lab_UT.didpuu0.countEnStens ),
            .ltout(\Lab_UT.didpuu0.countEnStens_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpstens.q_esr_ctle_3_LC_8_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpstens.q_esr_ctle_3_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpstens.q_esr_ctle_3_LC_8_7_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \Lab_UT.didpuu0.didpstens.q_esr_ctle_3_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12243),
            .in3(N__15919),
            .lcout(\Lab_UT.didpuu0.didpstens.countEnStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_0_LC_8_7_6 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_0_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpsones.q_0_LC_8_7_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_0_LC_8_7_6  (
            .in0(N__15691),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13307),
            .lcout(Lab_UT_di_Sones_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13519),
            .ce(),
            .sr(N__15885));
    defparam \uu2.un1_segment4_2_am_1_LC_8_7_7 .C_ON=1'b0;
    defparam \uu2.un1_segment4_2_am_1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_2_am_1_LC_8_7_7 .LUT_INIT=16'b0010010100000100;
    LogicCell40 \uu2.un1_segment4_2_am_1_LC_8_7_7  (
            .in0(N__14734),
            .in1(N__17237),
            .in2(N__14672),
            .in3(N__15689),
            .lcout(\uu2.un1_segment4_2_amZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNO_0_6_LC_8_8_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNO_0_6_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNO_0_6_LC_8_8_0 .LUT_INIT=16'b1011111011111010;
    LogicCell40 \uu2.w_addr_displaying_RNO_0_6_LC_8_8_0  (
            .in0(N__12338),
            .in1(N__12324),
            .in2(N__12225),
            .in3(N__13918),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_4_0_i_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_6_LC_8_8_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_LC_8_8_1 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_6_LC_8_8_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \uu2.w_addr_displaying_6_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__12212),
            .in2(N__12234),
            .in3(N__16057),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_6C_net ),
            .ce(),
            .sr(N__15849));
    defparam \uu2.w_addr_displaying_RNIKFL01_6_LC_8_8_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIKFL01_6_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIKFL01_6_LC_8_8_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uu2.w_addr_displaying_RNIKFL01_6_LC_8_8_2  (
            .in0(N__12523),
            .in1(N__12181),
            .in2(_gnd_net_),
            .in3(N__13781),
            .lcout(\uu2.g0_i_o4_0_a8_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_8_LC_8_8_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_LC_8_8_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_8_LC_8_8_3  (
            .in0(N__12534),
            .in1(N__16056),
            .in2(N__15309),
            .in3(N__15346),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_6C_net ),
            .ce(),
            .sr(N__15849));
    defparam \uu2.w_addr_displaying_fast_RNO_0_6_LC_8_8_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNO_0_6_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNO_0_6_LC_8_8_4 .LUT_INIT=16'b1011111011111010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNO_0_6_LC_8_8_4  (
            .in0(N__12337),
            .in1(N__12323),
            .in2(N__14573),
            .in3(N__13917),
            .lcout(\uu2.w_addr_displaying_4_0_i_fast_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIHKAF2_8_LC_8_8_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIHKAF2_8_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIHKAF2_8_LC_8_8_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIHKAF2_8_LC_8_8_5  (
            .in0(N__15301),
            .in1(N__12524),
            .in2(_gnd_net_),
            .in3(N__15345),
            .lcout(\uu2.un15_w_data_displaying ),
            .ltout(\uu2.un15_w_data_displaying_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIMF2HD_8_LC_8_8_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIMF2HD_8_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIMF2HD_8_LC_8_8_6 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \uu2.w_addr_displaying_RNIMF2HD_8_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12486),
            .in3(N__12426),
            .lcout(\uu2.un21_w_addr_displaying_i ),
            .ltout(\uu2.un21_w_addr_displaying_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_7_LC_8_8_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_LC_8_8_7 .LUT_INIT=16'b1100110001101100;
    LogicCell40 \uu2.w_addr_displaying_7_LC_8_8_7  (
            .in0(N__13919),
            .in1(N__16251),
            .in2(N__12345),
            .in3(N__14012),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_6C_net ),
            .ce(),
            .sr(N__15849));
    defparam \uu2.w_addr_displaying_6_rep1_LC_8_9_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_rep1_LC_8_9_0 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_6_rep1_LC_8_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.w_addr_displaying_6_rep1_LC_8_9_0  (
            .in0(N__16045),
            .in1(N__12252),
            .in2(_gnd_net_),
            .in3(N__16414),
            .lcout(\uu2.w_addr_displaying_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_6_rep1C_net ),
            .ce(),
            .sr(N__15853));
    defparam \uu2.w_addr_displaying_6_rep1_RNO_0_LC_8_9_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_rep1_RNO_0_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_6_rep1_RNO_0_LC_8_9_1 .LUT_INIT=16'b1111011011111010;
    LogicCell40 \uu2.w_addr_displaying_6_rep1_RNO_0_LC_8_9_1  (
            .in0(N__16413),
            .in1(N__13914),
            .in2(N__12342),
            .in3(N__12316),
            .lcout(\uu2.w_addr_displaying_4_0_i_rep1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_5_rep1_RNI3HMT_LC_8_9_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_rep1_RNI3HMT_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_5_rep1_RNI3HMT_LC_8_9_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uu2.w_addr_displaying_5_rep1_RNI3HMT_LC_8_9_2  (
            .in0(N__16409),
            .in1(N__16459),
            .in2(N__15456),
            .in3(N__15531),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_5_rep1_RNI3HMTZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_5_rep1_RNIMFM34_LC_8_9_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_rep1_RNIMFM34_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_5_rep1_RNIMFM34_LC_8_9_3 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \uu2.w_addr_displaying_5_rep1_RNIMFM34_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__13638),
            .in2(N__12246),
            .in3(N__14019),
            .lcout(\uu2.un1_segment3_m5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_5_LC_8_9_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_5_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_5_LC_8_9_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.w_addr_displaying_fast_5_LC_8_9_4  (
            .in0(N__13915),
            .in1(_gnd_net_),
            .in2(N__16091),
            .in3(N__14502),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_6_rep1C_net ),
            .ce(),
            .sr(N__15853));
    defparam \uu2.w_addr_displaying_fast_RNID5QH_5_LC_8_9_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNID5QH_5_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNID5QH_5_LC_8_9_5 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \uu2.w_addr_displaying_fast_RNID5QH_5_LC_8_9_5  (
            .in0(N__14500),
            .in1(N__14557),
            .in2(_gnd_net_),
            .in3(N__13822),
            .lcout(\uu2.w_addr_displaying_fast_RNID5QHZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI6N2K_5_LC_8_9_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI6N2K_5_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI6N2K_5_LC_8_9_6 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI6N2K_5_LC_8_9_6  (
            .in0(N__14558),
            .in1(N__14501),
            .in2(N__13843),
            .in3(N__15532),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_fast_RNI6N2KZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI76AF1_2_LC_8_9_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI76AF1_2_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI76AF1_2_LC_8_9_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI76AF1_2_LC_8_9_7  (
            .in0(N__12681),
            .in1(_gnd_net_),
            .in2(N__12675),
            .in3(N__12672),
            .lcout(\uu2.un1_segment4_sn_N_39_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI2VHC_4_LC_8_10_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI2VHC_4_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI2VHC_4_LC_8_10_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI2VHC_4_LC_8_10_0  (
            .in0(N__12986),
            .in1(N__13069),
            .in2(N__15247),
            .in3(N__14234),
            .lcout(\uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4 ),
            .ltout(\uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNILB202_4_LC_8_10_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNILB202_4_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNILB202_4_LC_8_10_1 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \uu2.w_addr_displaying_RNILB202_4_LC_8_10_1  (
            .in0(N__13756),
            .in1(N__13680),
            .in2(N__12648),
            .in3(N__14454),
            .lcout(\uu2.w_addr_displaying_RNILB202Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_rep1_RNIR94U_LC_8_10_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_RNIR94U_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_2_rep1_RNIR94U_LC_8_10_2 .LUT_INIT=16'b1010001010001010;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_RNIR94U_LC_8_10_2  (
            .in0(N__14453),
            .in1(N__15452),
            .in2(N__15546),
            .in3(N__16347),
            .lcout(\uu2.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep2_RNI75VM_LC_8_10_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep2_RNI75VM_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_4_rep2_RNI75VM_LC_8_10_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uu2.w_addr_displaying_4_rep2_RNI75VM_LC_8_10_3  (
            .in0(N__13828),
            .in1(N__15426),
            .in2(N__14889),
            .in3(N__15533),
            .lcout(\uu2.w_addr_displaying_4_rep2_RNI75VMZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_rep1_RNI4RA21_LC_8_10_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_RNI4RA21_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_2_rep1_RNI4RA21_LC_8_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_RNI4RA21_LC_8_10_4  (
            .in0(N__15425),
            .in1(N__13827),
            .in2(N__16364),
            .in3(N__14866),
            .lcout(\uu2.un1_w_addr_displaying_inv_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_3_LC_8_10_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_3_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_3_LC_8_10_5 .LUT_INIT=16'b0011110011001100;
    LogicCell40 \uu2.w_addr_displaying_fast_3_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__13077),
            .in2(N__15490),
            .in3(N__16090),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_3C_net ),
            .ce(),
            .sr(N__15855));
    defparam \uu2.w_addr_displaying_fast_RNIN0TS_4_LC_8_10_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIN0TS_4_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIN0TS_4_LC_8_10_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIN0TS_4_LC_8_10_6  (
            .in0(N__12985),
            .in1(N__14288),
            .in2(N__13082),
            .in3(N__16346),
            .lcout(\uu2.w_addr_displaying_fast_RNIN0TSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNILHHC_0_LC_8_10_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNILHHC_0_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNILHHC_0_LC_8_10_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNILHHC_0_LC_8_10_7  (
            .in0(N__13070),
            .in1(N__12987),
            .in2(N__12963),
            .in3(N__15945),
            .lcout(\uu2.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_1_LC_8_11_0 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_1_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpsones.q_1_LC_8_11_0 .LUT_INIT=16'b0100011001001100;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_1_LC_8_11_0  (
            .in0(N__13321),
            .in1(N__17210),
            .in2(N__12918),
            .in3(N__15714),
            .lcout(Lab_UT_di_Sones_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13493),
            .ce(),
            .sr(N__15888));
    defparam \Lab_UT.didpuu0.didpsones.q_2_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_2_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpsones.q_2_LC_8_11_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_2_LC_8_11_1  (
            .in0(N__15715),
            .in1(N__13322),
            .in2(N__17238),
            .in3(N__14720),
            .lcout(Lab_UT_di_Sones_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13493),
            .ce(),
            .sr(N__15888));
    defparam \Lab_UT.didpuu0.didpsones.q_3_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_3_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpsones.q_3_LC_8_11_3 .LUT_INIT=16'b1110111011000100;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_3_LC_8_11_3  (
            .in0(N__13323),
            .in1(N__14619),
            .in2(N__12891),
            .in3(N__12873),
            .lcout(Lab_UT_di_Sones_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13493),
            .ce(),
            .sr(N__15888));
    defparam \uu2.segment1_m_2_0_LC_8_11_4 .C_ON=1'b0;
    defparam \uu2.segment1_m_2_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \uu2.segment1_m_2_0_LC_8_11_4 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \uu2.segment1_m_2_0_LC_8_11_4  (
            .in0(N__14719),
            .in1(N__17209),
            .in2(N__14637),
            .in3(N__15713),
            .lcout(),
            .ltout(\uu2.segment1_m_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_7_rep1_RNIPUSD1_LC_8_11_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_rep1_RNIPUSD1_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_7_rep1_RNIPUSD1_LC_8_11_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \uu2.w_addr_displaying_7_rep1_RNIPUSD1_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12846),
            .in3(N__14896),
            .lcout(),
            .ltout(\uu2.segment1_m_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIBOM74_3_LC_8_11_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIBOM74_3_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIBOM74_3_LC_8_11_6 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \uu2.w_addr_displaying_RNIBOM74_3_LC_8_11_6  (
            .in0(N__15367),
            .in1(N__13278),
            .in2(N__12843),
            .in3(N__12836),
            .lcout(),
            .ltout(\uu2.un1_segment1_iv_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_rep1_RNI2NR6D_LC_8_11_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_RNI2NR6D_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_0_rep1_RNI2NR6D_LC_8_11_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_RNI2NR6D_LC_8_11_7  (
            .in0(N__14319),
            .in1(N__12741),
            .in2(N__12735),
            .in3(N__16209),
            .lcout(\uu2.un1_segment1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpstens.q_esr_2_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpstens.q_esr_2_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpstens.q_esr_2_LC_8_12_1 .LUT_INIT=16'b0110011011000100;
    LogicCell40 \Lab_UT.didpuu0.didpstens.q_esr_2_LC_8_12_1  (
            .in0(N__15640),
            .in1(N__14160),
            .in2(N__14090),
            .in3(N__17329),
            .lcout(Lab_UT_di_Stens_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13490),
            .ce(N__13119),
            .sr(N__15891));
    defparam \Lab_UT.didpuu0.didpstens.q_esr_3_LC_8_12_3 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpstens.q_esr_3_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpstens.q_esr_3_LC_8_12_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \Lab_UT.didpuu0.didpstens.q_esr_3_LC_8_12_3  (
            .in0(N__15641),
            .in1(N__14161),
            .in2(N__14091),
            .in3(N__17330),
            .lcout(Lab_UT_di_Stens_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13490),
            .ce(N__13119),
            .sr(N__15891));
    defparam \uu2.un1_segment4_3_bm_LC_8_12_4 .C_ON=1'b0;
    defparam \uu2.un1_segment4_3_bm_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_3_bm_LC_8_12_4 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \uu2.un1_segment4_3_bm_LC_8_12_4  (
            .in0(N__14158),
            .in1(N__17327),
            .in2(N__14088),
            .in3(N__15638),
            .lcout(\uu2.un1_segment4_3_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment4_3_am_LC_8_12_5 .C_ON=1'b0;
    defparam \uu2.un1_segment4_3_am_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment4_3_am_LC_8_12_5 .LUT_INIT=16'b0001101110110111;
    LogicCell40 \uu2.un1_segment4_3_am_LC_8_12_5  (
            .in0(N__15639),
            .in1(N__14159),
            .in2(N__14089),
            .in3(N__17328),
            .lcout(),
            .ltout(\uu2.un1_segment4_3_amZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_rep1_RNI8N8R6_LC_8_12_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_RNI8N8R6_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_0_rep1_RNI8N8R6_LC_8_12_6 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_RNI8N8R6_LC_8_12_6  (
            .in0(N__14306),
            .in1(N__13107),
            .in2(N__13101),
            .in3(N__13098),
            .lcout(),
            .ltout(\uu2.N_289_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIFU9M8_8_LC_8_12_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIFU9M8_8_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIFU9M8_8_LC_8_12_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIFU9M8_8_LC_8_12_7  (
            .in0(N__15561),
            .in1(_gnd_net_),
            .in2(N__13092),
            .in3(N__15195),
            .lcout(\uu2.w_addr_displaying_fast_RNIFU9M8Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIBHTT_3_LC_8_13_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIBHTT_3_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIBHTT_3_LC_8_13_0 .LUT_INIT=16'b1001010110101001;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIBHTT_3_LC_8_13_0  (
            .in0(N__16363),
            .in1(N__13081),
            .in2(N__15002),
            .in3(N__14826),
            .lcout(\uu2.N_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep1_RNIAVDB_0_LC_8_13_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep1_RNIAVDB_0_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_4_rep1_RNIAVDB_0_LC_8_13_1 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \uu2.w_addr_displaying_4_rep1_RNIAVDB_0_LC_8_13_1  (
            .in0(N__15450),
            .in1(_gnd_net_),
            .in2(N__14831),
            .in3(N__14906),
            .lcout(\uu2.w_addr_displaying_4_rep1_RNIAVDBZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIKFIE_6_LC_8_13_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIKFIE_6_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIKFIE_6_LC_8_13_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIKFIE_6_LC_8_13_2  (
            .in0(N__15547),
            .in1(N__15451),
            .in2(N__14907),
            .in3(N__14574),
            .lcout(\uu2.w_addr_displaying_fast_RNIKFIEZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMU_0_LC_8_13_3 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMU_0_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMU_0_LC_8_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMU_0_LC_8_13_3  (
            .in0(N__14071),
            .in1(N__14650),
            .in2(_gnd_net_),
            .in3(N__17111),
            .lcout(),
            .ltout(\Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMUZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIRNGO1_1_LC_8_13_4 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIRNGO1_1_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIRNGO1_1_LC_8_13_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNIRNGO1_1_LC_8_13_4  (
            .in0(N__13251),
            .in1(_gnd_net_),
            .in2(N__13266),
            .in3(N__17164),
            .lcout(led_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI67CI_0_LC_8_13_5 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI67CI_0_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI67CI_0_LC_8_13_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNI67CI_0_LC_8_13_5  (
            .in0(N__17110),
            .in1(N__16741),
            .in2(_gnd_net_),
            .in3(N__15099),
            .lcout(\Lab_UT.didpuu0.ledDisp00.selLed_RNI67CIZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec1.un11_segmentUQ_1_0_a2_LC_8_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dec1.un11_segmentUQ_1_0_a2_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec1.un11_segmentUQ_1_0_a2_LC_8_13_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dec1.un11_segmentUQ_1_0_a2_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__14167),
            .in2(_gnd_net_),
            .in3(N__14070),
            .lcout(\Lab_UT.un11_segmentUQ_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpmones.q_esr_RNIF7VF1_3_LC_8_14_0 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmones.q_esr_RNIF7VF1_3_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpmones.q_esr_RNIF7VF1_3_LC_8_14_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.didpuu0.didpmones.q_esr_RNIF7VF1_3_LC_8_14_0  (
            .in0(N__16930),
            .in1(N__16841),
            .in2(N__16782),
            .in3(N__16658),
            .lcout(),
            .ltout(\Lab_UT.didpuu0.countEnMtens_0_a4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpstens.q_RNIJUV53_1_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpstens.q_RNIJUV53_1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpstens.q_RNIJUV53_1_LC_8_14_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.didpuu0.didpstens.q_RNIJUV53_1_LC_8_14_1  (
            .in0(N__13229),
            .in1(N__17331),
            .in2(N__13218),
            .in3(N__15642),
            .lcout(\Lab_UT.didpuu0.countEnMtens_0_a4_1 ),
            .ltout(\Lab_UT.didpuu0.countEnMtens_0_a4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpstens.q_RNI4BA55_1_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpstens.q_RNI4BA55_1_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpstens.q_RNI4BA55_1_LC_8_14_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.didpuu0.didpstens.q_RNI4BA55_1_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13191),
            .in3(N__13188),
            .lcout(\Lab_UT.didpuu0.countEnMtens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpmones.q_2_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmones.q_2_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpmones.q_2_LC_8_14_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \Lab_UT.didpuu0.didpmones.q_2_LC_8_14_3  (
            .in0(N__16659),
            .in1(N__13656),
            .in2(N__16865),
            .in3(N__16931),
            .lcout(Lab_UT_di_Mones_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13485),
            .ce(),
            .sr(N__15894));
    defparam \uu2.segment3_m_3_1_LC_8_14_4 .C_ON=1'b0;
    defparam \uu2.segment3_m_3_1_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \uu2.segment3_m_3_1_LC_8_14_4 .LUT_INIT=16'b0011110101010111;
    LogicCell40 \uu2.segment3_m_3_1_LC_8_14_4  (
            .in0(N__16928),
            .in1(N__16840),
            .in2(N__16781),
            .in3(N__16657),
            .lcout(\uu2.segment3_m_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpmones.q_1_LC_8_14_5 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmones.q_1_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpmones.q_1_LC_8_14_5 .LUT_INIT=16'b0011010011110000;
    LogicCell40 \Lab_UT.didpuu0.didpmones.q_1_LC_8_14_5  (
            .in0(N__13125),
            .in1(N__16668),
            .in2(N__16866),
            .in3(N__13655),
            .lcout(Lab_UT_di_Mones_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13485),
            .ce(),
            .sr(N__15894));
    defparam \Lab_UT.didpuu0.didpmones.q_0_LC_8_14_6 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpmones.q_0_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpmones.q_0_LC_8_14_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.didpuu0.didpmones.q_0_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__13654),
            .in2(_gnd_net_),
            .in3(N__16660),
            .lcout(Lab_UT_di_Mones_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13485),
            .ce(),
            .sr(N__15894));
    defparam \uu2.un1_segment3_m5_bm_LC_8_14_7 .C_ON=1'b0;
    defparam \uu2.un1_segment3_m5_bm_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment3_m5_bm_LC_8_14_7 .LUT_INIT=16'b0101111010110101;
    LogicCell40 \uu2.un1_segment3_m5_bm_LC_8_14_7  (
            .in0(N__16656),
            .in1(N__16767),
            .in2(N__16864),
            .in3(N__16929),
            .lcout(\uu2.un1_segment3_m5_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_LC_9_5_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_0_LC_9_5_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_0_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__13622),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13539),
            .ce(N__13578),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.sec_clkD_LC_9_7_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.sec_clkD_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.secuu0.sec_clkD_LC_9_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.secuu0.sec_clkD_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16542),
            .lcout(\Lab_UT.sec_clkD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13526),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.clkSecStrb_LC_9_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.clkSecStrb_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.clkSecStrb_LC_9_7_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.didpuu0.clkSecStrb_LC_9_7_1  (
            .in0(N__16541),
            .in1(N__13334),
            .in2(_gnd_net_),
            .in3(N__16577),
            .lcout(\Lab_UT.didpuu0.clkSecStrbZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.segment2_m_2_5_LC_9_7_4 .C_ON=1'b0;
    defparam \uu2.segment2_m_2_5_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.segment2_m_2_5_LC_9_7_4 .LUT_INIT=16'b1101001011111011;
    LogicCell40 \uu2.segment2_m_2_5_LC_9_7_4  (
            .in0(N__14187),
            .in1(N__17299),
            .in2(N__14110),
            .in3(N__15610),
            .lcout(\uu2.segment2_m_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec1.segmentUQ_4_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dec1.segmentUQ_4_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec1.segmentUQ_4_LC_9_8_0 .LUT_INIT=16'b1111010111010001;
    LogicCell40 \Lab_UT.dec1.segmentUQ_4_LC_9_8_0  (
            .in0(N__15628),
            .in1(N__14190),
            .in2(N__14112),
            .in3(N__17317),
            .lcout(),
            .ltout(L3_segment2_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep1_RNIBG883_LC_9_8_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep1_RNIBG883_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_4_rep1_RNIBG883_LC_9_8_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \uu2.w_addr_displaying_4_rep1_RNIBG883_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__13293),
            .in2(N__13281),
            .in3(N__14791),
            .lcout(\uu2.un1_segment3_m0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.segment2_m_1_6_LC_9_8_2 .C_ON=1'b0;
    defparam \uu2.segment2_m_1_6_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.segment2_m_1_6_LC_9_8_2 .LUT_INIT=16'b1111011110111100;
    LogicCell40 \uu2.segment2_m_1_6_LC_9_8_2  (
            .in0(N__15627),
            .in1(N__14189),
            .in2(N__14111),
            .in3(N__17318),
            .lcout(\uu2.segment2_m_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_segment3_m5_am_LC_9_8_3 .C_ON=1'b0;
    defparam \uu2.un1_segment3_m5_am_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_segment3_m5_am_LC_9_8_3 .LUT_INIT=16'b0110011010111101;
    LogicCell40 \uu2.un1_segment3_m5_am_LC_9_8_3  (
            .in0(N__14188),
            .in1(N__17316),
            .in2(N__14113),
            .in3(N__15626),
            .lcout(\uu2.un1_segment3_m5_amZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep1_LC_9_8_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep1_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_rep1_LC_9_8_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.w_addr_displaying_4_rep1_LC_9_8_4  (
            .in0(N__14792),
            .in1(N__15305),
            .in2(_gnd_net_),
            .in3(N__16054),
            .lcout(\uu2.w_addr_displaying_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4_rep1C_net ),
            .ce(),
            .sr(N__15851));
    defparam \uu2.w_addr_displaying_fast_RNILLSO_7_LC_9_8_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNILLSO_7_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNILLSO_7_LC_9_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNILLSO_7_LC_9_8_5  (
            .in0(N__16458),
            .in1(N__14222),
            .in2(N__16417),
            .in3(N__14790),
            .lcout(\uu2.Z_decfrac106_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_5_rep1_LC_9_8_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_rep1_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_rep1_LC_9_8_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.w_addr_displaying_5_rep1_LC_9_8_6  (
            .in0(N__16463),
            .in1(N__13925),
            .in2(_gnd_net_),
            .in3(N__16055),
            .lcout(\uu2.w_addr_displaying_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4_rep1C_net ),
            .ce(),
            .sr(N__15851));
    defparam \uu2.w_addr_displaying_fast_7_LC_9_8_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_7_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_7_LC_9_8_7 .LUT_INIT=16'b1101111100100000;
    LogicCell40 \uu2.w_addr_displaying_fast_7_LC_9_8_7  (
            .in0(N__16053),
            .in1(N__14011),
            .in2(N__13929),
            .in3(N__14223),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4_rep1C_net ),
            .ce(),
            .sr(N__15851));
    defparam \uu2.w_addr_displaying_4_rep1_RNI65VM_LC_9_9_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep1_RNI65VM_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_4_rep1_RNI65VM_LC_9_9_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uu2.w_addr_displaying_4_rep1_RNI65VM_LC_9_9_0  (
            .in0(N__14820),
            .in1(N__15441),
            .in2(N__13857),
            .in3(N__14890),
            .lcout(\uu2.un1_w_addr_displaying_35_0 ),
            .ltout(\uu2.un1_w_addr_displaying_35_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIPHFA2_4_LC_9_9_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIPHFA2_4_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIPHFA2_4_LC_9_9_1 .LUT_INIT=16'b1111111111110010;
    LogicCell40 \uu2.w_addr_displaying_RNIPHFA2_4_LC_9_9_1  (
            .in0(N__14461),
            .in1(N__13779),
            .in2(N__13683),
            .in3(N__13679),
            .lcout(\uu2.N_813_0 ),
            .ltout(\uu2.N_813_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_9_9_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_9_9_2 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_58_LC_9_9_2  (
            .in0(N__16595),
            .in1(N__14415),
            .in2(N__13668),
            .in3(N__14369),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep1_RNIAVDB_LC_9_9_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep1_RNIAVDB_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_4_rep1_RNIAVDB_LC_9_9_3 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \uu2.w_addr_displaying_4_rep1_RNIAVDB_LC_9_9_3  (
            .in0(N__14891),
            .in1(N__14821),
            .in2(_gnd_net_),
            .in3(N__15442),
            .lcout(\uu2.un1_segment3_m4_s_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec0.segmentUQ_3_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dec0.segmentUQ_3_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec0.segmentUQ_3_LC_9_9_4 .LUT_INIT=16'b0110011010111101;
    LogicCell40 \Lab_UT.dec0.segmentUQ_3_LC_9_9_4  (
            .in0(N__14749),
            .in1(N__17239),
            .in2(N__14679),
            .in3(N__15725),
            .lcout(),
            .ltout(L3_segment1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIQD7R4_5_LC_9_9_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIQD7R4_5_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIQD7R4_5_LC_9_9_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIQD7R4_5_LC_9_9_5  (
            .in0(N__14580),
            .in1(N__14572),
            .in2(N__14514),
            .in3(N__14503),
            .lcout(\uu2.w_addr_displaying_fast_RNIQD7R4Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIL396_8_LC_9_9_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIL396_8_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIL396_8_LC_9_9_6 .LUT_INIT=16'b0000001100000011;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIL396_8_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__14221),
            .in2(N__15240),
            .in3(_gnd_net_),
            .lcout(\uu2.N_315_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_9_9_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_9_9_7 .LUT_INIT=16'b1101110111110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_59_LC_9_9_7  (
            .in0(N__14416),
            .in1(N__16596),
            .in2(N__14384),
            .in3(N__14346),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_rep1_RNIUV0B3_LC_9_10_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_RNIUV0B3_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_0_rep1_RNIUV0B3_LC_9_10_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_RNIUV0B3_LC_9_10_0  (
            .in0(N__16252),
            .in1(N__14286),
            .in2(N__14331),
            .in3(N__16491),
            .lcout(\uu2.segment2_m_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_rep1_LC_9_10_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_rep1_LC_9_10_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_LC_9_10_1  (
            .in0(N__14287),
            .in1(_gnd_net_),
            .in2(N__16095),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displaying_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0_rep1C_net ),
            .ce(),
            .sr(N__15856));
    defparam \uu2.w_addr_displaying_4_rep2_RNI4S6J_LC_9_10_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep2_RNI4S6J_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_4_rep2_RNI4S6J_LC_9_10_2 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \uu2.w_addr_displaying_4_rep2_RNI4S6J_LC_9_10_2  (
            .in0(N__15420),
            .in1(N__14284),
            .in2(_gnd_net_),
            .in3(N__15526),
            .lcout(\uu2.w_addr_displaying_4_rep2_RNI4S6JZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIEDBM_7_LC_9_10_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIEDBM_7_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIEDBM_7_LC_9_10_3 .LUT_INIT=16'b0010010000000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIEDBM_7_LC_9_10_3  (
            .in0(N__14285),
            .in1(N__15421),
            .in2(N__15545),
            .in3(N__14233),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_fast_RNIEDBMZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNITRMC1_8_LC_9_10_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNITRMC1_8_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNITRMC1_8_LC_9_10_4 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNITRMC1_8_LC_9_10_4  (
            .in0(N__15235),
            .in1(N__15570),
            .in2(N__15564),
            .in3(_gnd_net_),
            .lcout(\uu2.un1_segment4_sn_N_38_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep2_LC_9_10_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep2_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_rep2_LC_9_10_5 .LUT_INIT=16'b0110101001101010;
    LogicCell40 \uu2.w_addr_displaying_4_rep2_LC_9_10_5  (
            .in0(N__15530),
            .in1(N__15307),
            .in2(N__16096),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displaying_4_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0_rep1C_net ),
            .ce(),
            .sr(N__15856));
    defparam \uu2.w_addr_displaying_3_rep1_LC_9_10_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_rep1_LC_9_10_6 .LUT_INIT=16'b0011110011110000;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__15491),
            .in2(N__15449),
            .in3(N__16065),
            .lcout(\uu2.w_addr_displaying_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0_rep1C_net ),
            .ce(),
            .sr(N__15856));
    defparam \uu2.w_addr_displaying_fast_8_LC_9_10_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_8_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_8_LC_9_10_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_displaying_fast_8_LC_9_10_7  (
            .in0(N__16066),
            .in1(N__15236),
            .in2(N__15368),
            .in3(N__15308),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0_rep1C_net ),
            .ce(),
            .sr(N__15856));
    defparam \Lab_UT.dec3.segmentUQ_2_LC_9_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dec3.segmentUQ_2_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec3.segmentUQ_2_LC_9_11_0 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \Lab_UT.dec3.segmentUQ_2_LC_9_11_0  (
            .in0(N__15182),
            .in1(N__17050),
            .in2(N__15100),
            .in3(N__17443),
            .lcout(),
            .ltout(L3_segment4_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_rep1_RNIABAE_LC_9_11_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_RNIABAE_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_2_rep1_RNIABAE_LC_9_11_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_RNIABAE_LC_9_11_1  (
            .in0(N__16344),
            .in1(_gnd_net_),
            .in2(N__15198),
            .in3(N__15009),
            .lcout(\uu2.N_280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dec3.segmentUQ_4_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dec3.segmentUQ_4_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dec3.segmentUQ_4_LC_9_11_2 .LUT_INIT=16'b1110000011111101;
    LogicCell40 \Lab_UT.dec3.segmentUQ_4_LC_9_11_2  (
            .in0(N__15183),
            .in1(N__17049),
            .in2(N__15101),
            .in3(N__17442),
            .lcout(L3_segment4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_rep1_LC_9_11_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_rep1_LC_9_11_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_LC_9_11_3  (
            .in0(N__16345),
            .in1(N__16136),
            .in2(N__16097),
            .in3(N__15003),
            .lcout(\uu2.w_addr_displaying_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__15858));
    defparam \uu2.w_addr_displaying_5_rep1_RNI9Q311_0_LC_9_11_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_rep1_RNI9Q311_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_5_rep1_RNI9Q311_0_LC_9_11_4 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \uu2.w_addr_displaying_5_rep1_RNI9Q311_0_LC_9_11_4  (
            .in0(N__16465),
            .in1(N__16416),
            .in2(_gnd_net_),
            .in3(N__16342),
            .lcout(\uu2.un1_w_addr_displaying_46_1 ),
            .ltout(\uu2.un1_w_addr_displaying_46_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI8U3D2_0_LC_9_11_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8U3D2_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8U3D2_0_LC_9_11_5 .LUT_INIT=16'b0000001111001111;
    LogicCell40 \uu2.w_addr_displaying_RNI8U3D2_0_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__16135),
            .in2(N__16485),
            .in3(N__16311),
            .lcout(\uu2.w_addr_displaying_RNI8U3D2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_5_rep1_RNI9Q311_LC_9_11_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_rep1_RNI9Q311_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_5_rep1_RNI9Q311_LC_9_11_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \uu2.w_addr_displaying_5_rep1_RNI9Q311_LC_9_11_6  (
            .in0(N__16464),
            .in1(N__16415),
            .in2(_gnd_net_),
            .in3(N__16343),
            .lcout(\uu2.un1_w_addr_displaying_38_1 ),
            .ltout(\uu2.un1_w_addr_displaying_38_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIBSR63_7_LC_9_11_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIBSR63_7_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIBSR63_7_LC_9_11_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIBSR63_7_LC_9_11_7  (
            .in0(N__16305),
            .in1(N__16134),
            .in2(N__16293),
            .in3(N__16253),
            .lcout(\uu2.segment3_m_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_LC_9_12_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_9_12_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_displaying_0_LC_9_12_0  (
            .in0(N__16094),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16152),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0C_net ),
            .ce(),
            .sr(N__15859));
    defparam \uu2.w_addr_displaying_fast_0_LC_9_12_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_0_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_0_LC_9_12_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_fast_0_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__16093),
            .in2(_gnd_net_),
            .in3(N__15943),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0C_net ),
            .ce(),
            .sr(N__15859));
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_9_13_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_9_13_0 .LUT_INIT=16'b1001111111101101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_60_LC_9_13_0  (
            .in0(N__16938),
            .in1(N__16855),
            .in2(N__16681),
            .in3(N__16780),
            .lcout(\uu2.mem0.N_2160_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11_0_LC_9_13_2 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11_0_LC_9_13_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11_0_LC_9_13_2  (
            .in0(N__15735),
            .in1(N__17112),
            .in2(_gnd_net_),
            .in3(N__15654),
            .lcout(),
            .ltout(\Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNITQOS1_1_LC_9_13_3 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNITQOS1_1_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNITQOS1_1_LC_9_13_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNITQOS1_1_LC_9_13_3  (
            .in0(N__17166),
            .in1(_gnd_net_),
            .in2(N__17466),
            .in3(N__17349),
            .lcout(led_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNINURJ_0_LC_9_13_4 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNINURJ_0_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNINURJ_0_LC_9_13_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNINURJ_0_LC_9_13_4  (
            .in0(N__17451),
            .in1(N__16669),
            .in2(_gnd_net_),
            .in3(N__17114),
            .lcout(\Lab_UT.didpuu0.ledDisp00.selLed_RNINURJZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11_0_LC_9_13_5 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11_0_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11_0_LC_9_13_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11_0_LC_9_13_5  (
            .in0(N__17113),
            .in1(N__17343),
            .in2(_gnd_net_),
            .in3(N__17254),
            .lcout(),
            .ltout(\Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI1VOS1_1_LC_9_13_6 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI1VOS1_1_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNI1VOS1_1_LC_9_13_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNI1VOS1_1_LC_9_13_6  (
            .in0(N__16977),
            .in1(_gnd_net_),
            .in2(N__17169),
            .in3(N__17165),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJ_0_LC_9_13_7 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJ_0_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJ_0_LC_9_13_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJ_0_LC_9_13_7  (
            .in0(N__17115),
            .in1(_gnd_net_),
            .in2(N__16873),
            .in3(N__17062),
            .lcout(\Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.g0_i_0_LC_9_14_7 .C_ON=1'b0;
    defparam \uu2.g0_i_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \uu2.g0_i_0_LC_9_14_7 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \uu2.g0_i_0_LC_9_14_7  (
            .in0(N__16932),
            .in1(N__16848),
            .in2(N__16783),
            .in3(N__16661),
            .lcout(\uu2.N_2160_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.o_oneSecPluse_LC_11_9_0 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.o_oneSecPluse_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.o_oneSecPluse_LC_11_9_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didpuu0.o_oneSecPluse_LC_11_9_0  (
            .in0(N__16581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16548),
            .lcout(led_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // latticehx1k

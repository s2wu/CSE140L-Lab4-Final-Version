-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Feb 25 2020 07:08:25

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__13611\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13392\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal clk_in_c : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \resetGen.rst_isoZ0\ : std_logic;
signal \Lab_UT.secuu0.un131_ci_3_cascade_\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \Lab_UT.secuu0.un197_ci_9_cascade_\ : std_logic;
signal \Lab_UT.secuu0.un230_ci_1_cascade_\ : std_logic;
signal \Lab_UT.secuu0.l_precountZ0Z_0\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_4\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_14_cascade_\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_0_8\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_0_8_cascade_\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_14\ : std_logic;
signal \Lab_UT.secuu0.un197_ci_9\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_12\ : std_logic;
signal \Lab_UT.secuu0.un208_ci_0\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_13\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_10\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_8\ : std_logic;
signal \uu2.mem0.w_addr_8\ : std_logic;
signal \uu2.mem0.w_addr_1\ : std_logic;
signal \uu2.mem0.w_addr_2\ : std_logic;
signal \uu2.mem0.w_addr_5\ : std_logic;
signal \uu2.mem0.w_data_4\ : std_logic;
signal \uu2.mem0.w_addr_3\ : std_logic;
signal \uu2.mem0.g0_0_a3_3_cascade_\ : std_logic;
signal \uu2.mem0.w_data_1\ : std_logic;
signal \uu2.mem0.g1_0_6_cascade_\ : std_logic;
signal \uu2.mem0.N_4_i\ : std_logic;
signal \uu2.mem0.w_addr_6\ : std_logic;
signal \uu2.mem0.N_14_0\ : std_logic;
signal \uu2.vbuf_raddr.un459_ci_0_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \uu2.vbuf_raddr.un437_ci_3\ : std_logic;
signal \uu2.un306_ci_cascade_\ : std_logic;
signal \uu2.un339_ci_0\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal \uu2.un415_ci_0\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu2.un3_r_clk_en_6_cascade_\ : std_logic;
signal \uu2_un3_r_clk_en_0_cascade_\ : std_logic;
signal \uu2.vbuf_tx_data_rdy\ : std_logic;
signal \uu2.un3_r_clk_en_0_0\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal \uu2.un3_r_clk_en_7\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \uu2.un372_ci_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_10\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.vbuf_count.un372_ci_8_1\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \uu2.vbuf_count.un372_ci_8_1_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uu2.un306_ci\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \Lab_UT.secuu0.l_precountZ0Z_2\ : std_logic;
signal \Lab_UT.secuu0.l_precountZ0Z_1\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_5\ : std_logic;
signal \Lab_UT.secuu0.l_precountZ0Z_3\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_15\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_11_cascade_\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_13\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_16_cascade_\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_18\ : std_logic;
signal \Lab_UT.secuu0.delay_lineZ0Z_1\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_0_cascade_\ : std_logic;
signal \Lab_UT.secuu0.delay_lineZ0Z_0\ : std_logic;
signal \Lab_UT.secuu0.un11_l_count_i\ : std_logic;
signal \Lab_UT.secuu0.un186_ci_0\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_11\ : std_logic;
signal \Lab_UT.secuu0.un241_ci_2\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_16\ : std_logic;
signal \Lab_UT.secuu0.un263_ci_cascade_\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_18\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_9\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_17\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_12\ : std_logic;
signal \Lab_UT.secuu0.un87_ci\ : std_logic;
signal \Lab_UT.secuu0.un87_ci_cascade_\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_3\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_2\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_0\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_1\ : std_logic;
signal \Lab_UT.secuu0.un109_ci_cascade_\ : std_logic;
signal \Lab_UT.secuu0.un153_ci\ : std_logic;
signal \Lab_UT.secuu0.un131_ci_3\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_6\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_0\ : std_logic;
signal \Lab_UT.secuu0.un142_ci_0\ : std_logic;
signal \Lab_UT.secuu0.un109_ci\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_7\ : std_logic;
signal \Lab_UT.secuu0.un11_l_count_i_g\ : std_logic;
signal \resetGen.N_104_cascade_\ : std_logic;
signal \resetGen.N_84\ : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \resetGen.N_86\ : std_logic;
signal \resetGen.N_104\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \resetGen.N_86_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_4\ : std_logic;
signal \uu2.mem0.g2_1_0_0_cascade_\ : std_logic;
signal \uu2.mem0.g0_2_1\ : std_logic;
signal \uu2.mem0.g0_i_a2_3_cascade_\ : std_logic;
signal \uu2.mem0.w_data_displaying_2_0_0\ : std_logic;
signal \uu2.mem0.g1_0_5\ : std_logic;
signal \uu2.mem0.N_10_0_0\ : std_logic;
signal \uu2.mem0.g1_2\ : std_logic;
signal \uu2.mem0.g1_1_sx\ : std_logic;
signal \uu2.mem0.g1_0\ : std_logic;
signal \uu2.mem0.g0_i_5\ : std_logic;
signal \uu2.mem0.g0_i_6_1_0\ : std_logic;
signal \uu2.mem0.N_19_cascade_\ : std_logic;
signal \uu2.mem0.g0_i_6\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_53\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \uu2.mem0.g0_0_a3_0\ : std_logic;
signal \buart.Z_rx.startbit_cascade_\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_rx.ser_clk_cascade_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \uu2.vbuf_tx_data_rdy_0\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \uu2.mem0.w_data_7\ : std_logic;
signal \buart.Z_rx.ser_clk\ : std_logic;
signal \buart.Z_rx.N_103_cascade_\ : std_logic;
signal \resetGen.un3_reset_count_i_a3Z0Z_7\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_4\ : std_logic;
signal \N_87_cascade_\ : std_logic;
signal \buart.Z_rx.N_91\ : std_logic;
signal \buart.Z_rx.N_91_cascade_\ : std_logic;
signal \buart.Z_rx.N_29_0_i_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.N_29_0_i_2_cascade_\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_rx.bitcounte_0_i_2\ : std_logic;
signal \uu2.Z_decfrac105_7_3_cascade_\ : std_logic;
signal \uu2.mem0.w_data_6\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_17_cascade_\ : std_logic;
signal \uu2.mem0.w_data_5\ : std_logic;
signal \uu2.Z_decfrac105_7_3\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_\ : std_logic;
signal \uu2.mem0.w_data_0\ : std_logic;
signal \INVuu2.w_addr_displaying_5C_net\ : std_logic;
signal \uu2.mem0.w_data_2\ : std_logic;
signal \uu2.un1_w_user_cr_0_0\ : std_logic;
signal \latticehx1k_pll_inst_PLLOUTCORE_i\ : std_logic;
signal \uu2.un1_w_user_cr_0_0_cascade_\ : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_34_cascade_\ : std_logic;
signal \uu2.mem0.un1_segment3_m6_0_0_0_0_cascade_\ : std_logic;
signal \uu2.mem0.w_data_3\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_35\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_21\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_22\ : std_logic;
signal \uu2.mem0.g0_i_a2_4\ : std_logic;
signal \uu2.mem0.N_8_tz_0_0_1\ : std_logic;
signal \led_c_0_4_cascade_\ : std_logic;
signal \uu2.mem0.g1_0_0_0\ : std_logic;
signal \uu2.mem0.g0_i_5_1_0\ : std_logic;
signal \uu2.mem0.g2_0\ : std_logic;
signal \uu2.w_addr_displaying_4_rep1_8_cascade_\ : std_logic;
signal \uu2.N_42_0_0_cascade_\ : std_logic;
signal \uu2.N_1482_0_0\ : std_logic;
signal \INVuu2.w_addr_displaying_8_rep1C_net\ : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal \uu2.o_adder_vbuf_w_addr_user_3_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.w_addr_userZ1Z_1\ : std_logic;
signal \INVuu2.w_addr_user_2C_net\ : std_logic;
signal \uu2.o_adder_vbuf_w_addr_user_7_cascade_\ : std_logic;
signal \uu2.mem0.w_addr_7\ : std_logic;
signal \uu2.vbuf_w_addr_user.un459_ci_0_cascade_\ : std_logic;
signal \uu2.o_adder_vbuf_w_addr_user_8_cascade_\ : std_logic;
signal \INVuu2.w_addr_user_7C_net\ : std_logic;
signal \uu2.un437_ci_3\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \uu2.un2_w_addr_user_4_cascade_\ : std_logic;
signal \uu2.un2_w_addr_user_5\ : std_logic;
signal \uu2.un448_ci_5_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \uu2.un415_ci\ : std_logic;
signal \INVuu2.w_addr_user_5C_net\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \uu2.mem0.w_addr_4\ : std_logic;
signal \uu2.mem0.g0_8_0_cascade_\ : std_logic;
signal \uu2.mem0.w_data_ns_1_1_0_3_cascade_\ : std_logic;
signal \uu2.Z_decfrac106\ : std_logic;
signal \uu2.mem0.w_data_ns_1_0_0_1_3\ : std_logic;
signal \uu2.g0_1_0_0_1_cascade_\ : std_logic;
signal \uu2.g0_1_0_0\ : std_logic;
signal \INVuu2.w_addr_displaying_5_rep1C_net\ : std_logic;
signal \uu2.g0_1_a5_0_0\ : std_logic;
signal \uu2.g0_1_a5_1_0\ : std_logic;
signal \uu2.g1_1\ : std_logic;
signal \INVuu2.w_addr_displaying_2_rep1C_net\ : std_logic;
signal \uu2.w_addr_displaying_8_repZ0Z1\ : std_logic;
signal \uu2.g1_0_1_cascade_\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_50_cascade_\ : std_logic;
signal \uu2.g1_0_1\ : std_logic;
signal \uu2.mem0.g0_0\ : std_logic;
signal \uu2.w_addr_displaying_7_repZ0Z1\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_\ : std_logic;
signal \uu2.mem0.g1\ : std_logic;
signal \uu2.N_10\ : std_logic;
signal \uu2.mem0.g1_1_1\ : std_logic;
signal \INVuu2.w_addr_displaying_0_rep1C_net\ : std_logic;
signal \uu2.w_addr_displaying_0_repZ0Z1\ : std_logic;
signal \uu2.mem0.N_10_0\ : std_logic;
signal \uu2.w_addr_displaying_4_rep1_3_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_1_repZ0Z1\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_2\ : std_logic;
signal \uu2.mem0.un1_segment4_0_i_i_1\ : std_logic;
signal \INVuu2.w_addr_displaying_3_rep1C_net\ : std_logic;
signal \uu2.mem0.un1_segment4_0_i_i_a5_0_0\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.q13_0_cascade_\ : std_logic;
signal \uu2.g0_3Z0Z_0\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \INVuu2.w_addr_user_0C_net\ : std_logic;
signal \uu2.w_addr_user_2Z0Z_1_cascade_\ : std_logic;
signal \uu2.w_addr_userZ2Z_1_cascade_\ : std_logic;
signal \uu2.w_addr_user_RNIT1MGDZ0Z_4\ : std_logic;
signal \uu2.w_addr_user_1_0\ : std_logic;
signal \Lab_UT.dictrluu0.dek.det_NZ0Z_5_cascade_\ : std_logic;
signal \uu2.mem0.N_1476_0_0_0\ : std_logic;
signal \Lab_UT.dspStr.cnt11_1\ : std_logic;
signal \uu2.w_m5_i_a3Z0Z_2\ : std_logic;
signal \Lab_UT.dictrluu0.dek.det_NZ0Z_4\ : std_logic;
signal \uu2.un1_w_user_lf_0_0Z0Z_0_cascade_\ : std_logic;
signal \uu2.un1_w_user_lf_2\ : std_logic;
signal \uu2.un2_w_addr_user\ : std_logic;
signal \uu2.un1_w_user_lf_2_cascade_\ : std_logic;
signal \uu2.un27_N_6_mux_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \uu2.w_addr_user_RNILDNK6Z0Z_4_cascade_\ : std_logic;
signal \uu2.un27_w_addr_user_i\ : std_logic;
signal \uu2.un1_w_user_lf_5_a0Z0Z_5_cascade_\ : std_logic;
signal \uu2.un1_w_user_lf_5_aZ0Z0\ : std_logic;
signal \Lab_UT_dspStr_cnt_1_rep1\ : std_logic;
signal \Lab_UT_dspStr_un36_dOut\ : std_logic;
signal \Lab_UT_dspStr_un36_dOut_cascade_\ : std_logic;
signal \uu2.un27_N_6_mux_cascade_\ : std_logic;
signal \uu2.un27_w_addr_user_iZ0Z_1\ : std_logic;
signal \Lab_UT_dspStr_cnt_3_rep1\ : std_logic;
signal \Lab_UT_dspStr_cnt_2_rep1\ : std_logic;
signal \L3_tx_data_0\ : std_logic;
signal \L3_tx_data_0_cascade_\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_1\ : std_logic;
signal \uu2.w_addr_displaying_RNIQKOV8Z0Z_8_cascade_\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal \uu2.un21_w_addr_displaying_i_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_6C_net\ : std_logic;
signal \uu2.mem0.g0_i_a11_1_0\ : std_logic;
signal \uu2.w_addr_displaying_4_repZ0Z1\ : std_logic;
signal \uu2.mem0.g3_0_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_3_repZ0Z1\ : std_logic;
signal \uu2.mem0.un1_segment4_0_i_i_0_0\ : std_logic;
signal \uu2.mem0.g0_i_a11_3_1\ : std_logic;
signal \uu2.mem0.g0_i_a11_7_1_cascade_\ : std_logic;
signal \uu2.mem0.g0_i_5_1\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_0C_net\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_0\ : std_logic;
signal \uu2.w_addr_displaying_6_repZ0Z1\ : std_logic;
signal \uu2.w_addr_displaying_5_repZ0Z1\ : std_logic;
signal \uu2.mem0.bitmap_pmux_1_1_i_a5_1_0\ : std_logic;
signal \uu2.mem0.g1_1_0_cascade_\ : std_logic;
signal \uu2.Z_decfrac106_5\ : std_logic;
signal \uu2.mem0.g0_2_0\ : std_logic;
signal \uu2.mem0.bitmap_pmux_1_1_i_a5_2_3_1_0\ : std_logic;
signal \uu2.w_addr_displaying_2_repZ0Z1\ : std_logic;
signal \uu2.Z_decfrac105_7_2\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_1\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_1C_net\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_4\ : std_logic;
signal \uu2.mem0.Z_decfrac105_7_3_2\ : std_logic;
signal \uu2.w_addr_displaying_4_8_cascade_\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \uu2.un15_w_data_displaying\ : std_logic;
signal \uu2.un15_w_data_displaying_cascade_\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_7\ : std_logic;
signal \INVuu2.w_addr_displaying_8C_net\ : std_logic;
signal \uu2.un448_ci_5\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.un1_q_cry_0\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_2\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.un1_q_cry_1\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.un1_q_cry_2\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_0\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_1\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.q13_0\ : std_logic;
signal rst : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \buart.Z_tx.bitcount_RNO_0Z0Z_1\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_0\ : std_logic;
signal \buart.Z_tx.bitcount_RNO_0Z0Z_2\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_1\ : std_logic;
signal uu2_un3_r_clk_en_0 : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_2\ : std_logic;
signal \buart.Z_tx.bitcount_RNIM5O32Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart__tx_uart_busy_0_cascade_\ : std_logic;
signal \buart.Z_tx.bitcount_RNIL4O32Z0Z_1\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \buart__tx_uart_busy_0\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.un1_bitcount_axb_3\ : std_logic;
signal \Lab_UT.dspStr.cnt11_0_i\ : std_logic;
signal \Lab_UT.dspStr.cntZ0Z_0\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \Lab_UT.dspStr.un1_cnt_3_cry_0\ : std_logic;
signal \Lab_UT.dspStr.un1_cnt_3_cry_1\ : std_logic;
signal \Lab_UT.dspStr.un1_cnt_3_cry_2\ : std_logic;
signal \Lab_UT_dspStr_cnt_1\ : std_logic;
signal \buart__rx_bitcount_3\ : std_logic;
signal \buart__rx_bitcount_2\ : std_logic;
signal \N_87\ : std_logic;
signal \Lab_UT.rx_data_rdy\ : std_logic;
signal \buart__rx_bitcount_0\ : std_logic;
signal \resetGen.un3_reset_count_i_a3Z0Z_4\ : std_logic;
signal \Lab_UT_L3_tx_data_0_6\ : std_logic;
signal \Lab_UT_dspStr_cnt_2\ : std_logic;
signal \Lab_UT_dspStr_cnt_3\ : std_logic;
signal \Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9EZ0\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.un4_w_user_data_rdyZ0Z_0\ : std_logic;
signal \uu2.mem0.w_addr_0\ : std_logic;
signal \Lab_UT_L3_tx_data_0_5_cascade_\ : std_logic;
signal \Lab_UT_L3_tx_data_0_2_6\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_4\ : std_logic;
signal \Lab_UT_L3_tx_data_0_2_1\ : std_logic;
signal \Lab_UT_L3_tx_data_2_3\ : std_logic;
signal \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87EZ0\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \Lab_UT.dspStr.cnt_fastZ0Z_1\ : std_logic;
signal \Lab_UT.dspStr.cnt_fastZ0Z_3\ : std_logic;
signal \Lab_UT_L3_tx_data_0_4\ : std_logic;
signal \Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8EZ0\ : std_logic;
signal \Lab_UT.dspStr.cnt_fastZ0Z_2\ : std_logic;
signal \Lab_UT_rx_data_0\ : std_logic;
signal \Lab_UT_rx_data_1\ : std_logic;
signal \Lab_UT_rx_data_2\ : std_logic;
signal \Lab_UT_rx_data_3\ : std_logic;
signal \Lab_UT_rx_data_6\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_6\ : std_logic;
signal \uu2.mem0.N_13_0\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_3\ : std_logic;
signal \uu2.w_addr_displaying_4_3\ : std_logic;
signal \Lab_UT_rx_data_7\ : std_logic;
signal \Lab_UT_rx_data_5\ : std_logic;
signal \Lab_UT_rx_data_4\ : std_logic;
signal \uu2.un1_w_user_lf_5_a0Z0Z_4\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.un437_ci\ : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \Lab_UT.Lab3U00.bu_rx_data_rdy_0\ : std_logic;
signal \Lab_UT.sec_clkD\ : std_logic;
signal \Lab_UT.didpuu0.clkSecStrbZ0\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_3\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \uu2.w_addr_displaying_4_fast_3\ : std_logic;
signal \uu2.mem0.g0_i_a11_2_0\ : std_logic;
signal \uu2.un15_w_data_displaying_5\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_4\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_5\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.un21_w_addr_displaying_i\ : std_logic;
signal \uu2.w_addr_displaying_4_fast_8\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_8\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_5C_net\ : std_logic;
signal \resetGen_rst_iso_g\ : std_logic;
signal \resetGen.un3_reset_count_i_a3Z0Z_5\ : std_logic;
signal bu_rx_data_0 : std_logic;
signal bu_rx_data_1 : std_logic;
signal bu_rx_data_7 : std_logic;
signal bu_rx_data_6 : std_logic;
signal bu_rx_data_5 : std_logic;
signal bu_rx_data_4 : std_logic;
signal bu_rx_data_3 : std_logic;
signal bu_rx_data_2 : std_logic;
signal clk_g : std_logic;
signal \buart.Z_rx.N_57_i\ : std_logic;
signal \Lab_UT_di_Sones_0\ : std_logic;
signal led_c_0 : std_logic;
signal \Lab_UT_dicRun\ : std_logic;
signal \Lab_UT_l_oneSecPluse\ : std_logic;
signal led_c_4 : std_logic;
signal \Lab_UT_di_Sones_2\ : std_logic;
signal led_c_2 : std_logic;
signal \Lab_UT_di_Sones_3\ : std_logic;
signal led_c_3 : std_logic;
signal \Lab_UT.dicSelectLEDdisp\ : std_logic;
signal \Lab_UT_di_Sones_1\ : std_logic;
signal led_c_1 : std_logic;
signal \_gnd_net_\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__5510\&\N__5471\&\N__5495\&\N__5453\&\N__5423\&\N__5608\&\N__5639\&\N__5675\&\N__5579\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__5282\&\N__7898\&\N__5360\&\N__5252\&\N__7949\&\N__5237\&\N__5264\&\N__5273\&\N__11135\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&\N__7316\&'0'&\N__7355\&'0'&\N__7667\&'0'&\N__5243\&'0'&\N__7724\&'0'&\N__7634\&'0'&\N__5375\&'0'&\N__7646\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \latticehx1k_pll_inst_PLLOUTCORE_i\,
            REFERENCECLK => \N__5054\,
            RESETB => \N__8894\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => \N__5828\,
            RCLK => \N__13421\,
            RE => \N__5827\,
            WCLKE => \N__7588\,
            WCLK => \N__13420\,
            WE => \N__7592\
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13611\,
            DIN => \N__13610\,
            DOUT => \N__13609\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13611\,
            PADOUT => \N__13610\,
            PADIN => \N__13609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13076\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13602\,
            DIN => \N__13601\,
            DOUT => \N__13600\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13602\,
            PADOUT => \N__13601\,
            PADIN => \N__13600\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13593\,
            DIN => \N__13592\,
            DOUT => \N__13591\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13593\,
            PADOUT => \N__13592\,
            PADIN => \N__13591\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12818\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13584\,
            DIN => \N__13583\,
            DOUT => \N__13582\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13584\,
            PADOUT => \N__13583\,
            PADIN => \N__13582\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7187\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13575\,
            DIN => \N__13574\,
            DOUT => \N__13573\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13575\,
            PADOUT => \N__13574\,
            PADIN => \N__13573\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13566\,
            DIN => \N__13565\,
            DOUT => \N__13564\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13566\,
            PADOUT => \N__13565\,
            PADIN => \N__13564\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13010\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13557\,
            DIN => \N__13556\,
            DOUT => \N__13555\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13557\,
            PADOUT => \N__13556\,
            PADIN => \N__13555\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12932\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13548\,
            DIN => \N__13547\,
            DOUT => \N__13546\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13548\,
            PADOUT => \N__13547\,
            PADIN => \N__13546\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13178\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13539\,
            DIN => \N__13538\,
            DOUT => \N__13537\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__13539\,
            PADOUT => \N__13538\,
            PADIN => \N__13537\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__13415\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13530\,
            DIN => \N__13529\,
            DOUT => \N__13528\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13530\,
            PADOUT => \N__13529\,
            PADIN => \N__13528\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3253\ : InMux
    port map (
            O => \N__13511\,
            I => \N__13507\
        );

    \I__3252\ : InMux
    port map (
            O => \N__13510\,
            I => \N__13503\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__13507\,
            I => \N__13500\
        );

    \I__3250\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13497\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__13503\,
            I => \N__13492\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__13500\,
            I => \N__13492\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__13497\,
            I => bu_rx_data_4
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__13492\,
            I => bu_rx_data_4
        );

    \I__3245\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13483\
        );

    \I__3244\ : InMux
    port map (
            O => \N__13486\,
            I => \N__13480\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__13483\,
            I => \N__13474\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__13480\,
            I => \N__13474\
        );

    \I__3241\ : InMux
    port map (
            O => \N__13479\,
            I => \N__13471\
        );

    \I__3240\ : Span4Mux_v
    port map (
            O => \N__13474\,
            I => \N__13468\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__13471\,
            I => bu_rx_data_3
        );

    \I__3238\ : Odrv4
    port map (
            O => \N__13468\,
            I => bu_rx_data_3
        );

    \I__3237\ : InMux
    port map (
            O => \N__13463\,
            I => \N__13459\
        );

    \I__3236\ : InMux
    port map (
            O => \N__13462\,
            I => \N__13456\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__13459\,
            I => \N__13453\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__13456\,
            I => \N__13449\
        );

    \I__3233\ : Span4Mux_v
    port map (
            O => \N__13453\,
            I => \N__13446\
        );

    \I__3232\ : InMux
    port map (
            O => \N__13452\,
            I => \N__13443\
        );

    \I__3231\ : Span4Mux_v
    port map (
            O => \N__13449\,
            I => \N__13438\
        );

    \I__3230\ : Span4Mux_h
    port map (
            O => \N__13446\,
            I => \N__13438\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__13443\,
            I => bu_rx_data_2
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__13438\,
            I => bu_rx_data_2
        );

    \I__3227\ : ClkMux
    port map (
            O => \N__13433\,
            I => \N__13265\
        );

    \I__3226\ : ClkMux
    port map (
            O => \N__13432\,
            I => \N__13265\
        );

    \I__3225\ : ClkMux
    port map (
            O => \N__13431\,
            I => \N__13265\
        );

    \I__3224\ : ClkMux
    port map (
            O => \N__13430\,
            I => \N__13265\
        );

    \I__3223\ : ClkMux
    port map (
            O => \N__13429\,
            I => \N__13265\
        );

    \I__3222\ : ClkMux
    port map (
            O => \N__13428\,
            I => \N__13265\
        );

    \I__3221\ : ClkMux
    port map (
            O => \N__13427\,
            I => \N__13265\
        );

    \I__3220\ : ClkMux
    port map (
            O => \N__13426\,
            I => \N__13265\
        );

    \I__3219\ : ClkMux
    port map (
            O => \N__13425\,
            I => \N__13265\
        );

    \I__3218\ : ClkMux
    port map (
            O => \N__13424\,
            I => \N__13265\
        );

    \I__3217\ : ClkMux
    port map (
            O => \N__13423\,
            I => \N__13265\
        );

    \I__3216\ : ClkMux
    port map (
            O => \N__13422\,
            I => \N__13265\
        );

    \I__3215\ : ClkMux
    port map (
            O => \N__13421\,
            I => \N__13265\
        );

    \I__3214\ : ClkMux
    port map (
            O => \N__13420\,
            I => \N__13265\
        );

    \I__3213\ : ClkMux
    port map (
            O => \N__13419\,
            I => \N__13265\
        );

    \I__3212\ : ClkMux
    port map (
            O => \N__13418\,
            I => \N__13265\
        );

    \I__3211\ : ClkMux
    port map (
            O => \N__13417\,
            I => \N__13265\
        );

    \I__3210\ : ClkMux
    port map (
            O => \N__13416\,
            I => \N__13265\
        );

    \I__3209\ : ClkMux
    port map (
            O => \N__13415\,
            I => \N__13265\
        );

    \I__3208\ : ClkMux
    port map (
            O => \N__13414\,
            I => \N__13265\
        );

    \I__3207\ : ClkMux
    port map (
            O => \N__13413\,
            I => \N__13265\
        );

    \I__3206\ : ClkMux
    port map (
            O => \N__13412\,
            I => \N__13265\
        );

    \I__3205\ : ClkMux
    port map (
            O => \N__13411\,
            I => \N__13265\
        );

    \I__3204\ : ClkMux
    port map (
            O => \N__13410\,
            I => \N__13265\
        );

    \I__3203\ : ClkMux
    port map (
            O => \N__13409\,
            I => \N__13265\
        );

    \I__3202\ : ClkMux
    port map (
            O => \N__13408\,
            I => \N__13265\
        );

    \I__3201\ : ClkMux
    port map (
            O => \N__13407\,
            I => \N__13265\
        );

    \I__3200\ : ClkMux
    port map (
            O => \N__13406\,
            I => \N__13265\
        );

    \I__3199\ : ClkMux
    port map (
            O => \N__13405\,
            I => \N__13265\
        );

    \I__3198\ : ClkMux
    port map (
            O => \N__13404\,
            I => \N__13265\
        );

    \I__3197\ : ClkMux
    port map (
            O => \N__13403\,
            I => \N__13265\
        );

    \I__3196\ : ClkMux
    port map (
            O => \N__13402\,
            I => \N__13265\
        );

    \I__3195\ : ClkMux
    port map (
            O => \N__13401\,
            I => \N__13265\
        );

    \I__3194\ : ClkMux
    port map (
            O => \N__13400\,
            I => \N__13265\
        );

    \I__3193\ : ClkMux
    port map (
            O => \N__13399\,
            I => \N__13265\
        );

    \I__3192\ : ClkMux
    port map (
            O => \N__13398\,
            I => \N__13265\
        );

    \I__3191\ : ClkMux
    port map (
            O => \N__13397\,
            I => \N__13265\
        );

    \I__3190\ : ClkMux
    port map (
            O => \N__13396\,
            I => \N__13265\
        );

    \I__3189\ : ClkMux
    port map (
            O => \N__13395\,
            I => \N__13265\
        );

    \I__3188\ : ClkMux
    port map (
            O => \N__13394\,
            I => \N__13265\
        );

    \I__3187\ : ClkMux
    port map (
            O => \N__13393\,
            I => \N__13265\
        );

    \I__3186\ : ClkMux
    port map (
            O => \N__13392\,
            I => \N__13265\
        );

    \I__3185\ : ClkMux
    port map (
            O => \N__13391\,
            I => \N__13265\
        );

    \I__3184\ : ClkMux
    port map (
            O => \N__13390\,
            I => \N__13265\
        );

    \I__3183\ : ClkMux
    port map (
            O => \N__13389\,
            I => \N__13265\
        );

    \I__3182\ : ClkMux
    port map (
            O => \N__13388\,
            I => \N__13265\
        );

    \I__3181\ : ClkMux
    port map (
            O => \N__13387\,
            I => \N__13265\
        );

    \I__3180\ : ClkMux
    port map (
            O => \N__13386\,
            I => \N__13265\
        );

    \I__3179\ : ClkMux
    port map (
            O => \N__13385\,
            I => \N__13265\
        );

    \I__3178\ : ClkMux
    port map (
            O => \N__13384\,
            I => \N__13265\
        );

    \I__3177\ : ClkMux
    port map (
            O => \N__13383\,
            I => \N__13265\
        );

    \I__3176\ : ClkMux
    port map (
            O => \N__13382\,
            I => \N__13265\
        );

    \I__3175\ : ClkMux
    port map (
            O => \N__13381\,
            I => \N__13265\
        );

    \I__3174\ : ClkMux
    port map (
            O => \N__13380\,
            I => \N__13265\
        );

    \I__3173\ : ClkMux
    port map (
            O => \N__13379\,
            I => \N__13265\
        );

    \I__3172\ : ClkMux
    port map (
            O => \N__13378\,
            I => \N__13265\
        );

    \I__3171\ : GlobalMux
    port map (
            O => \N__13265\,
            I => \N__13262\
        );

    \I__3170\ : gio2CtrlBuf
    port map (
            O => \N__13262\,
            I => clk_g
        );

    \I__3169\ : CEMux
    port map (
            O => \N__13259\,
            I => \N__13256\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__13256\,
            I => \N__13252\
        );

    \I__3167\ : CEMux
    port map (
            O => \N__13255\,
            I => \N__13249\
        );

    \I__3166\ : Span4Mux_v
    port map (
            O => \N__13252\,
            I => \N__13246\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__13249\,
            I => \N__13243\
        );

    \I__3164\ : Span4Mux_s2_h
    port map (
            O => \N__13246\,
            I => \N__13240\
        );

    \I__3163\ : Span4Mux_v
    port map (
            O => \N__13243\,
            I => \N__13237\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__13240\,
            I => \buart.Z_rx.N_57_i\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__13237\,
            I => \buart.Z_rx.N_57_i\
        );

    \I__3160\ : InMux
    port map (
            O => \N__13232\,
            I => \N__13229\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__13229\,
            I => \N__13220\
        );

    \I__3158\ : InMux
    port map (
            O => \N__13228\,
            I => \N__13211\
        );

    \I__3157\ : InMux
    port map (
            O => \N__13227\,
            I => \N__13211\
        );

    \I__3156\ : InMux
    port map (
            O => \N__13226\,
            I => \N__13211\
        );

    \I__3155\ : InMux
    port map (
            O => \N__13225\,
            I => \N__13211\
        );

    \I__3154\ : InMux
    port map (
            O => \N__13224\,
            I => \N__13205\
        );

    \I__3153\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13202\
        );

    \I__3152\ : Span4Mux_v
    port map (
            O => \N__13220\,
            I => \N__13199\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__13211\,
            I => \N__13196\
        );

    \I__3150\ : InMux
    port map (
            O => \N__13210\,
            I => \N__13189\
        );

    \I__3149\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13189\
        );

    \I__3148\ : InMux
    port map (
            O => \N__13208\,
            I => \N__13189\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__13205\,
            I => \Lab_UT_di_Sones_0\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__13202\,
            I => \Lab_UT_di_Sones_0\
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__13199\,
            I => \Lab_UT_di_Sones_0\
        );

    \I__3144\ : Odrv12
    port map (
            O => \N__13196\,
            I => \Lab_UT_di_Sones_0\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__13189\,
            I => \Lab_UT_di_Sones_0\
        );

    \I__3142\ : IoInMux
    port map (
            O => \N__13178\,
            I => \N__13175\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__13175\,
            I => \N__13172\
        );

    \I__3140\ : Odrv12
    port map (
            O => \N__13172\,
            I => led_c_0
        );

    \I__3139\ : InMux
    port map (
            O => \N__13169\,
            I => \N__13165\
        );

    \I__3138\ : InMux
    port map (
            O => \N__13168\,
            I => \N__13162\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__13165\,
            I => \N__13155\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__13162\,
            I => \N__13155\
        );

    \I__3135\ : InMux
    port map (
            O => \N__13161\,
            I => \N__13150\
        );

    \I__3134\ : InMux
    port map (
            O => \N__13160\,
            I => \N__13150\
        );

    \I__3133\ : Odrv12
    port map (
            O => \N__13155\,
            I => \Lab_UT_dicRun\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__13150\,
            I => \Lab_UT_dicRun\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__13145\,
            I => \N__13141\
        );

    \I__3130\ : InMux
    port map (
            O => \N__13144\,
            I => \N__13137\
        );

    \I__3129\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13131\
        );

    \I__3128\ : InMux
    port map (
            O => \N__13140\,
            I => \N__13131\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__13137\,
            I => \N__13128\
        );

    \I__3126\ : InMux
    port map (
            O => \N__13136\,
            I => \N__13125\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__13131\,
            I => \N__13122\
        );

    \I__3124\ : Span4Mux_v
    port map (
            O => \N__13128\,
            I => \N__13118\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__13125\,
            I => \N__13114\
        );

    \I__3122\ : Span4Mux_h
    port map (
            O => \N__13122\,
            I => \N__13111\
        );

    \I__3121\ : InMux
    port map (
            O => \N__13121\,
            I => \N__13108\
        );

    \I__3120\ : Span4Mux_v
    port map (
            O => \N__13118\,
            I => \N__13104\
        );

    \I__3119\ : InMux
    port map (
            O => \N__13117\,
            I => \N__13101\
        );

    \I__3118\ : Span4Mux_v
    port map (
            O => \N__13114\,
            I => \N__13094\
        );

    \I__3117\ : Span4Mux_v
    port map (
            O => \N__13111\,
            I => \N__13094\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__13108\,
            I => \N__13094\
        );

    \I__3115\ : InMux
    port map (
            O => \N__13107\,
            I => \N__13091\
        );

    \I__3114\ : Sp12to4
    port map (
            O => \N__13104\,
            I => \N__13086\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__13101\,
            I => \N__13086\
        );

    \I__3112\ : Span4Mux_h
    port map (
            O => \N__13094\,
            I => \N__13083\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__13091\,
            I => \Lab_UT_l_oneSecPluse\
        );

    \I__3110\ : Odrv12
    port map (
            O => \N__13086\,
            I => \Lab_UT_l_oneSecPluse\
        );

    \I__3109\ : Odrv4
    port map (
            O => \N__13083\,
            I => \Lab_UT_l_oneSecPluse\
        );

    \I__3108\ : IoInMux
    port map (
            O => \N__13076\,
            I => \N__13073\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__13073\,
            I => \N__13070\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__13070\,
            I => led_c_4
        );

    \I__3105\ : InMux
    port map (
            O => \N__13067\,
            I => \N__13062\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__13066\,
            I => \N__13059\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__13065\,
            I => \N__13056\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__13062\,
            I => \N__13051\
        );

    \I__3101\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13044\
        );

    \I__3100\ : InMux
    port map (
            O => \N__13056\,
            I => \N__13044\
        );

    \I__3099\ : InMux
    port map (
            O => \N__13055\,
            I => \N__13044\
        );

    \I__3098\ : InMux
    port map (
            O => \N__13054\,
            I => \N__13041\
        );

    \I__3097\ : Span4Mux_v
    port map (
            O => \N__13051\,
            I => \N__13033\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__13044\,
            I => \N__13033\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__13041\,
            I => \N__13033\
        );

    \I__3094\ : InMux
    port map (
            O => \N__13040\,
            I => \N__13027\
        );

    \I__3093\ : Span4Mux_h
    port map (
            O => \N__13033\,
            I => \N__13024\
        );

    \I__3092\ : InMux
    port map (
            O => \N__13032\,
            I => \N__13017\
        );

    \I__3091\ : InMux
    port map (
            O => \N__13031\,
            I => \N__13017\
        );

    \I__3090\ : InMux
    port map (
            O => \N__13030\,
            I => \N__13017\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__13027\,
            I => \Lab_UT_di_Sones_2\
        );

    \I__3088\ : Odrv4
    port map (
            O => \N__13024\,
            I => \Lab_UT_di_Sones_2\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__13017\,
            I => \Lab_UT_di_Sones_2\
        );

    \I__3086\ : IoInMux
    port map (
            O => \N__13010\,
            I => \N__13007\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__13007\,
            I => \N__13004\
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__13004\,
            I => led_c_2
        );

    \I__3083\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12995\
        );

    \I__3082\ : CascadeMux
    port map (
            O => \N__13000\,
            I => \N__12992\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__12999\,
            I => \N__12988\
        );

    \I__3080\ : CascadeMux
    port map (
            O => \N__12998\,
            I => \N__12985\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__12995\,
            I => \N__12980\
        );

    \I__3078\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12976\
        );

    \I__3077\ : InMux
    port map (
            O => \N__12991\,
            I => \N__12967\
        );

    \I__3076\ : InMux
    port map (
            O => \N__12988\,
            I => \N__12967\
        );

    \I__3075\ : InMux
    port map (
            O => \N__12985\,
            I => \N__12967\
        );

    \I__3074\ : InMux
    port map (
            O => \N__12984\,
            I => \N__12967\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__12983\,
            I => \N__12963\
        );

    \I__3072\ : Span4Mux_h
    port map (
            O => \N__12980\,
            I => \N__12959\
        );

    \I__3071\ : InMux
    port map (
            O => \N__12979\,
            I => \N__12956\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__12976\,
            I => \N__12953\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__12967\,
            I => \N__12950\
        );

    \I__3068\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12943\
        );

    \I__3067\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12943\
        );

    \I__3066\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12943\
        );

    \I__3065\ : Odrv4
    port map (
            O => \N__12959\,
            I => \Lab_UT_di_Sones_3\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__12956\,
            I => \Lab_UT_di_Sones_3\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__12953\,
            I => \Lab_UT_di_Sones_3\
        );

    \I__3062\ : Odrv12
    port map (
            O => \N__12950\,
            I => \Lab_UT_di_Sones_3\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__12943\,
            I => \Lab_UT_di_Sones_3\
        );

    \I__3060\ : IoInMux
    port map (
            O => \N__12932\,
            I => \N__12929\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__12929\,
            I => \N__12926\
        );

    \I__3058\ : Odrv4
    port map (
            O => \N__12926\,
            I => led_c_3
        );

    \I__3057\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12920\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__12920\,
            I => \N__12916\
        );

    \I__3055\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12911\
        );

    \I__3054\ : Span4Mux_v
    port map (
            O => \N__12916\,
            I => \N__12908\
        );

    \I__3053\ : InMux
    port map (
            O => \N__12915\,
            I => \N__12903\
        );

    \I__3052\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12903\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__12911\,
            I => \N__12900\
        );

    \I__3050\ : Sp12to4
    port map (
            O => \N__12908\,
            I => \N__12895\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__12903\,
            I => \N__12895\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__12900\,
            I => \N__12892\
        );

    \I__3047\ : Span12Mux_s4_h
    port map (
            O => \N__12895\,
            I => \N__12889\
        );

    \I__3046\ : Span4Mux_v
    port map (
            O => \N__12892\,
            I => \N__12886\
        );

    \I__3045\ : Odrv12
    port map (
            O => \N__12889\,
            I => \Lab_UT.dicSelectLEDdisp\
        );

    \I__3044\ : Odrv4
    port map (
            O => \N__12886\,
            I => \Lab_UT.dicSelectLEDdisp\
        );

    \I__3043\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12877\
        );

    \I__3042\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12868\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__12877\,
            I => \N__12864\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__12876\,
            I => \N__12861\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__12875\,
            I => \N__12857\
        );

    \I__3038\ : InMux
    port map (
            O => \N__12874\,
            I => \N__12848\
        );

    \I__3037\ : InMux
    port map (
            O => \N__12873\,
            I => \N__12848\
        );

    \I__3036\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12848\
        );

    \I__3035\ : InMux
    port map (
            O => \N__12871\,
            I => \N__12848\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__12868\,
            I => \N__12845\
        );

    \I__3033\ : InMux
    port map (
            O => \N__12867\,
            I => \N__12842\
        );

    \I__3032\ : Span4Mux_s3_h
    port map (
            O => \N__12864\,
            I => \N__12839\
        );

    \I__3031\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12832\
        );

    \I__3030\ : InMux
    port map (
            O => \N__12860\,
            I => \N__12832\
        );

    \I__3029\ : InMux
    port map (
            O => \N__12857\,
            I => \N__12832\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__12848\,
            I => \N__12829\
        );

    \I__3027\ : Odrv12
    port map (
            O => \N__12845\,
            I => \Lab_UT_di_Sones_1\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__12842\,
            I => \Lab_UT_di_Sones_1\
        );

    \I__3025\ : Odrv4
    port map (
            O => \N__12839\,
            I => \Lab_UT_di_Sones_1\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__12832\,
            I => \Lab_UT_di_Sones_1\
        );

    \I__3023\ : Odrv12
    port map (
            O => \N__12829\,
            I => \Lab_UT_di_Sones_1\
        );

    \I__3022\ : IoInMux
    port map (
            O => \N__12818\,
            I => \N__12815\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__12815\,
            I => \N__12812\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__12812\,
            I => led_c_1
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__12809\,
            I => \N__12805\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__12808\,
            I => \N__12799\
        );

    \I__3017\ : InMux
    port map (
            O => \N__12805\,
            I => \N__12793\
        );

    \I__3016\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12788\
        );

    \I__3015\ : InMux
    port map (
            O => \N__12803\,
            I => \N__12784\
        );

    \I__3014\ : InMux
    port map (
            O => \N__12802\,
            I => \N__12777\
        );

    \I__3013\ : InMux
    port map (
            O => \N__12799\,
            I => \N__12777\
        );

    \I__3012\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12777\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__12797\,
            I => \N__12774\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__12796\,
            I => \N__12770\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__12793\,
            I => \N__12766\
        );

    \I__3008\ : InMux
    port map (
            O => \N__12792\,
            I => \N__12763\
        );

    \I__3007\ : InMux
    port map (
            O => \N__12791\,
            I => \N__12760\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__12788\,
            I => \N__12756\
        );

    \I__3005\ : InMux
    port map (
            O => \N__12787\,
            I => \N__12753\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__12784\,
            I => \N__12748\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__12777\,
            I => \N__12748\
        );

    \I__3002\ : InMux
    port map (
            O => \N__12774\,
            I => \N__12739\
        );

    \I__3001\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12739\
        );

    \I__3000\ : InMux
    port map (
            O => \N__12770\,
            I => \N__12739\
        );

    \I__2999\ : InMux
    port map (
            O => \N__12769\,
            I => \N__12739\
        );

    \I__2998\ : Span4Mux_h
    port map (
            O => \N__12766\,
            I => \N__12732\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__12763\,
            I => \N__12732\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__12760\,
            I => \N__12732\
        );

    \I__2995\ : InMux
    port map (
            O => \N__12759\,
            I => \N__12729\
        );

    \I__2994\ : Span12Mux_s8_v
    port map (
            O => \N__12756\,
            I => \N__12726\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__12753\,
            I => \N__12719\
        );

    \I__2992\ : Span4Mux_h
    port map (
            O => \N__12748\,
            I => \N__12719\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__12739\,
            I => \N__12719\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__12732\,
            I => \uu2.un15_w_data_displaying_5\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__12729\,
            I => \uu2.un15_w_data_displaying_5\
        );

    \I__2988\ : Odrv12
    port map (
            O => \N__12726\,
            I => \uu2.un15_w_data_displaying_5\
        );

    \I__2987\ : Odrv4
    port map (
            O => \N__12719\,
            I => \uu2.un15_w_data_displaying_5\
        );

    \I__2986\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12707\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__12707\,
            I => \N__12702\
        );

    \I__2984\ : InMux
    port map (
            O => \N__12706\,
            I => \N__12699\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__12705\,
            I => \N__12695\
        );

    \I__2982\ : Span4Mux_v
    port map (
            O => \N__12702\,
            I => \N__12687\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__12699\,
            I => \N__12687\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__12698\,
            I => \N__12678\
        );

    \I__2979\ : InMux
    port map (
            O => \N__12695\,
            I => \N__12672\
        );

    \I__2978\ : InMux
    port map (
            O => \N__12694\,
            I => \N__12669\
        );

    \I__2977\ : InMux
    port map (
            O => \N__12693\,
            I => \N__12664\
        );

    \I__2976\ : InMux
    port map (
            O => \N__12692\,
            I => \N__12664\
        );

    \I__2975\ : Span4Mux_h
    port map (
            O => \N__12687\,
            I => \N__12661\
        );

    \I__2974\ : InMux
    port map (
            O => \N__12686\,
            I => \N__12658\
        );

    \I__2973\ : InMux
    port map (
            O => \N__12685\,
            I => \N__12651\
        );

    \I__2972\ : InMux
    port map (
            O => \N__12684\,
            I => \N__12651\
        );

    \I__2971\ : InMux
    port map (
            O => \N__12683\,
            I => \N__12651\
        );

    \I__2970\ : InMux
    port map (
            O => \N__12682\,
            I => \N__12644\
        );

    \I__2969\ : InMux
    port map (
            O => \N__12681\,
            I => \N__12644\
        );

    \I__2968\ : InMux
    port map (
            O => \N__12678\,
            I => \N__12644\
        );

    \I__2967\ : InMux
    port map (
            O => \N__12677\,
            I => \N__12637\
        );

    \I__2966\ : InMux
    port map (
            O => \N__12676\,
            I => \N__12637\
        );

    \I__2965\ : InMux
    port map (
            O => \N__12675\,
            I => \N__12637\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__12672\,
            I => \N__12634\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__12669\,
            I => \N__12629\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__12664\,
            I => \N__12629\
        );

    \I__2961\ : Odrv4
    port map (
            O => \N__12661\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__12658\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__12651\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__12644\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__12637\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2956\ : Odrv12
    port map (
            O => \N__12634\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2955\ : Odrv4
    port map (
            O => \N__12629\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2954\ : InMux
    port map (
            O => \N__12614\,
            I => \N__12610\
        );

    \I__2953\ : InMux
    port map (
            O => \N__12613\,
            I => \N__12607\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__12610\,
            I => \uu2.w_addr_displaying_fastZ0Z_5\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__12607\,
            I => \uu2.w_addr_displaying_fastZ0Z_5\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__12602\,
            I => \N__12595\
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__12601\,
            I => \N__12592\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__12600\,
            I => \N__12587\
        );

    \I__2947\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12581\
        );

    \I__2946\ : InMux
    port map (
            O => \N__12598\,
            I => \N__12576\
        );

    \I__2945\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12576\
        );

    \I__2944\ : InMux
    port map (
            O => \N__12592\,
            I => \N__12567\
        );

    \I__2943\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12567\
        );

    \I__2942\ : InMux
    port map (
            O => \N__12590\,
            I => \N__12567\
        );

    \I__2941\ : InMux
    port map (
            O => \N__12587\,
            I => \N__12567\
        );

    \I__2940\ : InMux
    port map (
            O => \N__12586\,
            I => \N__12564\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__12585\,
            I => \N__12558\
        );

    \I__2938\ : InMux
    port map (
            O => \N__12584\,
            I => \N__12555\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__12581\,
            I => \N__12550\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__12576\,
            I => \N__12550\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__12567\,
            I => \N__12547\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__12564\,
            I => \N__12544\
        );

    \I__2933\ : InMux
    port map (
            O => \N__12563\,
            I => \N__12541\
        );

    \I__2932\ : InMux
    port map (
            O => \N__12562\,
            I => \N__12538\
        );

    \I__2931\ : InMux
    port map (
            O => \N__12561\,
            I => \N__12533\
        );

    \I__2930\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12533\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__12555\,
            I => \N__12530\
        );

    \I__2928\ : Span4Mux_v
    port map (
            O => \N__12550\,
            I => \N__12525\
        );

    \I__2927\ : Span4Mux_v
    port map (
            O => \N__12547\,
            I => \N__12525\
        );

    \I__2926\ : Span4Mux_h
    port map (
            O => \N__12544\,
            I => \N__12522\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__12541\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__12538\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__12533\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2922\ : Odrv12
    port map (
            O => \N__12530\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__12525\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2920\ : Odrv4
    port map (
            O => \N__12522\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__12509\,
            I => \N__12505\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__12508\,
            I => \N__12490\
        );

    \I__2917\ : InMux
    port map (
            O => \N__12505\,
            I => \N__12476\
        );

    \I__2916\ : InMux
    port map (
            O => \N__12504\,
            I => \N__12476\
        );

    \I__2915\ : InMux
    port map (
            O => \N__12503\,
            I => \N__12476\
        );

    \I__2914\ : InMux
    port map (
            O => \N__12502\,
            I => \N__12476\
        );

    \I__2913\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12469\
        );

    \I__2912\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12469\
        );

    \I__2911\ : InMux
    port map (
            O => \N__12499\,
            I => \N__12469\
        );

    \I__2910\ : InMux
    port map (
            O => \N__12498\,
            I => \N__12457\
        );

    \I__2909\ : InMux
    port map (
            O => \N__12497\,
            I => \N__12457\
        );

    \I__2908\ : InMux
    port map (
            O => \N__12496\,
            I => \N__12450\
        );

    \I__2907\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12450\
        );

    \I__2906\ : InMux
    port map (
            O => \N__12494\,
            I => \N__12450\
        );

    \I__2905\ : InMux
    port map (
            O => \N__12493\,
            I => \N__12447\
        );

    \I__2904\ : InMux
    port map (
            O => \N__12490\,
            I => \N__12442\
        );

    \I__2903\ : InMux
    port map (
            O => \N__12489\,
            I => \N__12442\
        );

    \I__2902\ : InMux
    port map (
            O => \N__12488\,
            I => \N__12433\
        );

    \I__2901\ : InMux
    port map (
            O => \N__12487\,
            I => \N__12433\
        );

    \I__2900\ : InMux
    port map (
            O => \N__12486\,
            I => \N__12433\
        );

    \I__2899\ : InMux
    port map (
            O => \N__12485\,
            I => \N__12433\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__12476\,
            I => \N__12428\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__12469\,
            I => \N__12428\
        );

    \I__2896\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12423\
        );

    \I__2895\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12423\
        );

    \I__2894\ : InMux
    port map (
            O => \N__12466\,
            I => \N__12420\
        );

    \I__2893\ : InMux
    port map (
            O => \N__12465\,
            I => \N__12417\
        );

    \I__2892\ : InMux
    port map (
            O => \N__12464\,
            I => \N__12410\
        );

    \I__2891\ : InMux
    port map (
            O => \N__12463\,
            I => \N__12410\
        );

    \I__2890\ : InMux
    port map (
            O => \N__12462\,
            I => \N__12410\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__12457\,
            I => \N__12407\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__12450\,
            I => \N__12404\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__12447\,
            I => \N__12401\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__12442\,
            I => \N__12394\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__12433\,
            I => \N__12394\
        );

    \I__2884\ : Span4Mux_h
    port map (
            O => \N__12428\,
            I => \N__12394\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__12423\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__12420\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__12417\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__12410\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2879\ : Odrv4
    port map (
            O => \N__12407\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__12404\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__12401\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__12394\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2875\ : InMux
    port map (
            O => \N__12377\,
            I => \N__12374\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__12374\,
            I => \uu2.w_addr_displaying_4_fast_8\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__12371\,
            I => \N__12367\
        );

    \I__2872\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12362\
        );

    \I__2871\ : InMux
    port map (
            O => \N__12367\,
            I => \N__12362\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__12362\,
            I => \N__12359\
        );

    \I__2869\ : Span4Mux_h
    port map (
            O => \N__12359\,
            I => \N__12352\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__12358\,
            I => \N__12349\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__12357\,
            I => \N__12346\
        );

    \I__2866\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12343\
        );

    \I__2865\ : InMux
    port map (
            O => \N__12355\,
            I => \N__12340\
        );

    \I__2864\ : Span4Mux_s3_h
    port map (
            O => \N__12352\,
            I => \N__12337\
        );

    \I__2863\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12332\
        );

    \I__2862\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12332\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__12343\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__12340\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__12337\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__12332\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__2857\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12318\
        );

    \I__2856\ : SRMux
    port map (
            O => \N__12322\,
            I => \N__12313\
        );

    \I__2855\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12313\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__12318\,
            I => \N__12295\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__12313\,
            I => \N__12292\
        );

    \I__2852\ : SRMux
    port map (
            O => \N__12312\,
            I => \N__12224\
        );

    \I__2851\ : SRMux
    port map (
            O => \N__12311\,
            I => \N__12224\
        );

    \I__2850\ : SRMux
    port map (
            O => \N__12310\,
            I => \N__12224\
        );

    \I__2849\ : SRMux
    port map (
            O => \N__12309\,
            I => \N__12224\
        );

    \I__2848\ : SRMux
    port map (
            O => \N__12308\,
            I => \N__12224\
        );

    \I__2847\ : SRMux
    port map (
            O => \N__12307\,
            I => \N__12224\
        );

    \I__2846\ : SRMux
    port map (
            O => \N__12306\,
            I => \N__12224\
        );

    \I__2845\ : SRMux
    port map (
            O => \N__12305\,
            I => \N__12224\
        );

    \I__2844\ : SRMux
    port map (
            O => \N__12304\,
            I => \N__12224\
        );

    \I__2843\ : SRMux
    port map (
            O => \N__12303\,
            I => \N__12224\
        );

    \I__2842\ : SRMux
    port map (
            O => \N__12302\,
            I => \N__12224\
        );

    \I__2841\ : SRMux
    port map (
            O => \N__12301\,
            I => \N__12224\
        );

    \I__2840\ : SRMux
    port map (
            O => \N__12300\,
            I => \N__12224\
        );

    \I__2839\ : SRMux
    port map (
            O => \N__12299\,
            I => \N__12224\
        );

    \I__2838\ : SRMux
    port map (
            O => \N__12298\,
            I => \N__12224\
        );

    \I__2837\ : Glb2LocalMux
    port map (
            O => \N__12295\,
            I => \N__12224\
        );

    \I__2836\ : Glb2LocalMux
    port map (
            O => \N__12292\,
            I => \N__12224\
        );

    \I__2835\ : SRMux
    port map (
            O => \N__12291\,
            I => \N__12224\
        );

    \I__2834\ : SRMux
    port map (
            O => \N__12290\,
            I => \N__12224\
        );

    \I__2833\ : SRMux
    port map (
            O => \N__12289\,
            I => \N__12224\
        );

    \I__2832\ : SRMux
    port map (
            O => \N__12288\,
            I => \N__12224\
        );

    \I__2831\ : SRMux
    port map (
            O => \N__12287\,
            I => \N__12224\
        );

    \I__2830\ : SRMux
    port map (
            O => \N__12286\,
            I => \N__12224\
        );

    \I__2829\ : SRMux
    port map (
            O => \N__12285\,
            I => \N__12224\
        );

    \I__2828\ : SRMux
    port map (
            O => \N__12284\,
            I => \N__12224\
        );

    \I__2827\ : SRMux
    port map (
            O => \N__12283\,
            I => \N__12224\
        );

    \I__2826\ : SRMux
    port map (
            O => \N__12282\,
            I => \N__12224\
        );

    \I__2825\ : SRMux
    port map (
            O => \N__12281\,
            I => \N__12224\
        );

    \I__2824\ : GlobalMux
    port map (
            O => \N__12224\,
            I => \N__12221\
        );

    \I__2823\ : gio2CtrlBuf
    port map (
            O => \N__12221\,
            I => \resetGen_rst_iso_g\
        );

    \I__2822\ : InMux
    port map (
            O => \N__12218\,
            I => \N__12215\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__12215\,
            I => \N__12212\
        );

    \I__2820\ : Span4Mux_h
    port map (
            O => \N__12212\,
            I => \N__12209\
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__12209\,
            I => \resetGen.un3_reset_count_i_a3Z0Z_5\
        );

    \I__2818\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12203\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__12203\,
            I => \N__12199\
        );

    \I__2816\ : InMux
    port map (
            O => \N__12202\,
            I => \N__12196\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__12199\,
            I => bu_rx_data_0
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__12196\,
            I => bu_rx_data_0
        );

    \I__2813\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12188\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__12188\,
            I => \N__12183\
        );

    \I__2811\ : InMux
    port map (
            O => \N__12187\,
            I => \N__12178\
        );

    \I__2810\ : InMux
    port map (
            O => \N__12186\,
            I => \N__12178\
        );

    \I__2809\ : Odrv4
    port map (
            O => \N__12183\,
            I => bu_rx_data_1
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__12178\,
            I => bu_rx_data_1
        );

    \I__2807\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12169\
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__12172\,
            I => \N__12165\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__12169\,
            I => \N__12162\
        );

    \I__2804\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12159\
        );

    \I__2803\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12156\
        );

    \I__2802\ : Span4Mux_s3_h
    port map (
            O => \N__12162\,
            I => \N__12151\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__12159\,
            I => \N__12151\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__12156\,
            I => \N__12148\
        );

    \I__2799\ : Span4Mux_v
    port map (
            O => \N__12151\,
            I => \N__12145\
        );

    \I__2798\ : Span4Mux_v
    port map (
            O => \N__12148\,
            I => \N__12142\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__12145\,
            I => bu_rx_data_7
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__12142\,
            I => bu_rx_data_7
        );

    \I__2795\ : InMux
    port map (
            O => \N__12137\,
            I => \N__12133\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__12136\,
            I => \N__12129\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__12133\,
            I => \N__12126\
        );

    \I__2792\ : InMux
    port map (
            O => \N__12132\,
            I => \N__12121\
        );

    \I__2791\ : InMux
    port map (
            O => \N__12129\,
            I => \N__12121\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__12126\,
            I => bu_rx_data_6
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__12121\,
            I => bu_rx_data_6
        );

    \I__2788\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12113\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__12113\,
            I => \N__12108\
        );

    \I__2786\ : InMux
    port map (
            O => \N__12112\,
            I => \N__12103\
        );

    \I__2785\ : InMux
    port map (
            O => \N__12111\,
            I => \N__12103\
        );

    \I__2784\ : Odrv12
    port map (
            O => \N__12108\,
            I => bu_rx_data_5
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__12103\,
            I => bu_rx_data_5
        );

    \I__2782\ : InMux
    port map (
            O => \N__12098\,
            I => \N__12094\
        );

    \I__2781\ : InMux
    port map (
            O => \N__12097\,
            I => \N__12091\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__12094\,
            I => \uu2.w_addr_displaying_fastZ0Z_6\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__12091\,
            I => \uu2.w_addr_displaying_fastZ0Z_6\
        );

    \I__2778\ : InMux
    port map (
            O => \N__12086\,
            I => \N__12083\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__12083\,
            I => \uu2.mem0.N_13_0\
        );

    \I__2776\ : InMux
    port map (
            O => \N__12080\,
            I => \N__12074\
        );

    \I__2775\ : InMux
    port map (
            O => \N__12079\,
            I => \N__12069\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__12078\,
            I => \N__12066\
        );

    \I__2773\ : InMux
    port map (
            O => \N__12077\,
            I => \N__12060\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__12074\,
            I => \N__12056\
        );

    \I__2771\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12051\
        );

    \I__2770\ : InMux
    port map (
            O => \N__12072\,
            I => \N__12051\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__12069\,
            I => \N__12046\
        );

    \I__2768\ : InMux
    port map (
            O => \N__12066\,
            I => \N__12043\
        );

    \I__2767\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12038\
        );

    \I__2766\ : InMux
    port map (
            O => \N__12064\,
            I => \N__12038\
        );

    \I__2765\ : InMux
    port map (
            O => \N__12063\,
            I => \N__12035\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__12060\,
            I => \N__12032\
        );

    \I__2763\ : InMux
    port map (
            O => \N__12059\,
            I => \N__12029\
        );

    \I__2762\ : Span4Mux_v
    port map (
            O => \N__12056\,
            I => \N__12024\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__12051\,
            I => \N__12024\
        );

    \I__2760\ : InMux
    port map (
            O => \N__12050\,
            I => \N__12019\
        );

    \I__2759\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12019\
        );

    \I__2758\ : Span4Mux_h
    port map (
            O => \N__12046\,
            I => \N__12012\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__12043\,
            I => \N__12012\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__12038\,
            I => \N__12012\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__12035\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2754\ : Odrv4
    port map (
            O => \N__12032\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__12029\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2752\ : Odrv4
    port map (
            O => \N__12024\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__12019\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2750\ : Odrv4
    port map (
            O => \N__12012\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2749\ : InMux
    port map (
            O => \N__11999\,
            I => \N__11996\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__11996\,
            I => \N__11993\
        );

    \I__2747\ : Span4Mux_v
    port map (
            O => \N__11993\,
            I => \N__11990\
        );

    \I__2746\ : Span4Mux_h
    port map (
            O => \N__11990\,
            I => \N__11987\
        );

    \I__2745\ : Odrv4
    port map (
            O => \N__11987\,
            I => \uu2.w_addr_displaying_4_3\
        );

    \I__2744\ : InMux
    port map (
            O => \N__11984\,
            I => \N__11979\
        );

    \I__2743\ : InMux
    port map (
            O => \N__11983\,
            I => \N__11974\
        );

    \I__2742\ : InMux
    port map (
            O => \N__11982\,
            I => \N__11974\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__11979\,
            I => \N__11971\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__11974\,
            I => \N__11968\
        );

    \I__2739\ : Span4Mux_h
    port map (
            O => \N__11971\,
            I => \N__11963\
        );

    \I__2738\ : Span4Mux_h
    port map (
            O => \N__11968\,
            I => \N__11960\
        );

    \I__2737\ : InMux
    port map (
            O => \N__11967\,
            I => \N__11957\
        );

    \I__2736\ : InMux
    port map (
            O => \N__11966\,
            I => \N__11954\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__11963\,
            I => \Lab_UT_rx_data_7\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__11960\,
            I => \Lab_UT_rx_data_7\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__11957\,
            I => \Lab_UT_rx_data_7\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__11954\,
            I => \Lab_UT_rx_data_7\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__11945\,
            I => \N__11941\
        );

    \I__2730\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11938\
        );

    \I__2729\ : InMux
    port map (
            O => \N__11941\,
            I => \N__11935\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__11938\,
            I => \N__11931\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__11935\,
            I => \N__11928\
        );

    \I__2726\ : InMux
    port map (
            O => \N__11934\,
            I => \N__11925\
        );

    \I__2725\ : Span4Mux_h
    port map (
            O => \N__11931\,
            I => \N__11919\
        );

    \I__2724\ : Span4Mux_h
    port map (
            O => \N__11928\,
            I => \N__11919\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__11925\,
            I => \N__11916\
        );

    \I__2722\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11913\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__11919\,
            I => \Lab_UT_rx_data_5\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__11916\,
            I => \Lab_UT_rx_data_5\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__11913\,
            I => \Lab_UT_rx_data_5\
        );

    \I__2718\ : InMux
    port map (
            O => \N__11906\,
            I => \N__11900\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11905\,
            I => \N__11900\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__11900\,
            I => \N__11895\
        );

    \I__2715\ : InMux
    port map (
            O => \N__11899\,
            I => \N__11892\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11898\,
            I => \N__11889\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__11895\,
            I => \Lab_UT_rx_data_4\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__11892\,
            I => \Lab_UT_rx_data_4\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__11889\,
            I => \Lab_UT_rx_data_4\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11879\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__11879\,
            I => \N__11876\
        );

    \I__2708\ : Odrv4
    port map (
            O => \N__11876\,
            I => \uu2.un1_w_user_lf_5_a0Z0Z_4\
        );

    \I__2707\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11869\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11866\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__11869\,
            I => \N__11860\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__11866\,
            I => \N__11857\
        );

    \I__2703\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11852\
        );

    \I__2702\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11852\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__11863\,
            I => \N__11849\
        );

    \I__2700\ : Span4Mux_v
    port map (
            O => \N__11860\,
            I => \N__11840\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__11857\,
            I => \N__11840\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__11852\,
            I => \N__11840\
        );

    \I__2697\ : InMux
    port map (
            O => \N__11849\,
            I => \N__11835\
        );

    \I__2696\ : InMux
    port map (
            O => \N__11848\,
            I => \N__11835\
        );

    \I__2695\ : InMux
    port map (
            O => \N__11847\,
            I => \N__11832\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__11840\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__11835\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__11832\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__11825\,
            I => \N__11822\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11822\,
            I => \N__11819\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__11819\,
            I => \N__11814\
        );

    \I__2688\ : InMux
    port map (
            O => \N__11818\,
            I => \N__11811\
        );

    \I__2687\ : InMux
    port map (
            O => \N__11817\,
            I => \N__11808\
        );

    \I__2686\ : Span4Mux_h
    port map (
            O => \N__11814\,
            I => \N__11803\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__11811\,
            I => \N__11803\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__11808\,
            I => \N__11800\
        );

    \I__2683\ : Odrv4
    port map (
            O => \N__11803\,
            I => \uu2.un437_ci\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__11800\,
            I => \uu2.un437_ci\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11791\
        );

    \I__2680\ : InMux
    port map (
            O => \N__11794\,
            I => \N__11788\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11791\,
            I => \N__11785\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__11788\,
            I => \N__11782\
        );

    \I__2677\ : Span4Mux_v
    port map (
            O => \N__11785\,
            I => \N__11778\
        );

    \I__2676\ : Span4Mux_h
    port map (
            O => \N__11782\,
            I => \N__11775\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11772\
        );

    \I__2674\ : Odrv4
    port map (
            O => \N__11778\,
            I => bu_rx_data_rdy
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__11775\,
            I => bu_rx_data_rdy
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__11772\,
            I => bu_rx_data_rdy
        );

    \I__2671\ : CEMux
    port map (
            O => \N__11765\,
            I => \N__11762\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__11762\,
            I => \N__11759\
        );

    \I__2669\ : Odrv12
    port map (
            O => \N__11759\,
            I => \Lab_UT.Lab3U00.bu_rx_data_rdy_0\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__11756\,
            I => \N__11752\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11749\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11752\,
            I => \N__11746\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__11749\,
            I => \N__11743\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11746\,
            I => \N__11740\
        );

    \I__2663\ : Span4Mux_v
    port map (
            O => \N__11743\,
            I => \N__11735\
        );

    \I__2662\ : Span4Mux_h
    port map (
            O => \N__11740\,
            I => \N__11735\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__11735\,
            I => \Lab_UT.sec_clkD\
        );

    \I__2660\ : InMux
    port map (
            O => \N__11732\,
            I => \N__11726\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11721\
        );

    \I__2658\ : InMux
    port map (
            O => \N__11730\,
            I => \N__11721\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__11729\,
            I => \N__11716\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__11726\,
            I => \N__11711\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__11721\,
            I => \N__11711\
        );

    \I__2654\ : InMux
    port map (
            O => \N__11720\,
            I => \N__11704\
        );

    \I__2653\ : InMux
    port map (
            O => \N__11719\,
            I => \N__11704\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11704\
        );

    \I__2651\ : Span4Mux_h
    port map (
            O => \N__11711\,
            I => \N__11699\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__11704\,
            I => \N__11699\
        );

    \I__2649\ : Odrv4
    port map (
            O => \N__11699\,
            I => \Lab_UT.didpuu0.clkSecStrbZ0\
        );

    \I__2648\ : InMux
    port map (
            O => \N__11696\,
            I => \N__11687\
        );

    \I__2647\ : InMux
    port map (
            O => \N__11695\,
            I => \N__11687\
        );

    \I__2646\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11684\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11678\
        );

    \I__2644\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11678\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__11687\,
            I => \N__11671\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__11684\,
            I => \N__11668\
        );

    \I__2641\ : InMux
    port map (
            O => \N__11683\,
            I => \N__11665\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__11678\,
            I => \N__11662\
        );

    \I__2639\ : InMux
    port map (
            O => \N__11677\,
            I => \N__11653\
        );

    \I__2638\ : InMux
    port map (
            O => \N__11676\,
            I => \N__11653\
        );

    \I__2637\ : InMux
    port map (
            O => \N__11675\,
            I => \N__11653\
        );

    \I__2636\ : InMux
    port map (
            O => \N__11674\,
            I => \N__11653\
        );

    \I__2635\ : Span4Mux_s3_h
    port map (
            O => \N__11671\,
            I => \N__11646\
        );

    \I__2634\ : Span4Mux_v
    port map (
            O => \N__11668\,
            I => \N__11646\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__11665\,
            I => \N__11646\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__11662\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__11653\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__11646\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__11639\,
            I => \N__11634\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__11638\,
            I => \N__11630\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__11637\,
            I => \N__11624\
        );

    \I__2626\ : InMux
    port map (
            O => \N__11634\,
            I => \N__11621\
        );

    \I__2625\ : InMux
    port map (
            O => \N__11633\,
            I => \N__11618\
        );

    \I__2624\ : InMux
    port map (
            O => \N__11630\,
            I => \N__11609\
        );

    \I__2623\ : InMux
    port map (
            O => \N__11629\,
            I => \N__11609\
        );

    \I__2622\ : InMux
    port map (
            O => \N__11628\,
            I => \N__11609\
        );

    \I__2621\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11609\
        );

    \I__2620\ : InMux
    port map (
            O => \N__11624\,
            I => \N__11606\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__11621\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__11618\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__11609\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__11606\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__11597\,
            I => \N__11593\
        );

    \I__2614\ : InMux
    port map (
            O => \N__11596\,
            I => \N__11587\
        );

    \I__2613\ : InMux
    port map (
            O => \N__11593\,
            I => \N__11583\
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__11592\,
            I => \N__11580\
        );

    \I__2611\ : InMux
    port map (
            O => \N__11591\,
            I => \N__11575\
        );

    \I__2610\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11575\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__11587\,
            I => \N__11572\
        );

    \I__2608\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11568\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__11583\,
            I => \N__11565\
        );

    \I__2606\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11561\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__11575\,
            I => \N__11558\
        );

    \I__2604\ : Span4Mux_h
    port map (
            O => \N__11572\,
            I => \N__11555\
        );

    \I__2603\ : InMux
    port map (
            O => \N__11571\,
            I => \N__11552\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__11568\,
            I => \N__11547\
        );

    \I__2601\ : Span4Mux_h
    port map (
            O => \N__11565\,
            I => \N__11547\
        );

    \I__2600\ : InMux
    port map (
            O => \N__11564\,
            I => \N__11544\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__11561\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__11558\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__11555\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__11552\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__11547\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__11544\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2593\ : InMux
    port map (
            O => \N__11531\,
            I => \N__11528\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__11528\,
            I => \N__11525\
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__11525\,
            I => \uu2.w_addr_displaying_4_fast_3\
        );

    \I__2590\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11519\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__11519\,
            I => \N__11516\
        );

    \I__2588\ : Odrv4
    port map (
            O => \N__11516\,
            I => \uu2.mem0.g0_i_a11_2_0\
        );

    \I__2587\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11510\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__11510\,
            I => \N__11506\
        );

    \I__2585\ : InMux
    port map (
            O => \N__11509\,
            I => \N__11503\
        );

    \I__2584\ : Sp12to4
    port map (
            O => \N__11506\,
            I => \N__11497\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__11503\,
            I => \N__11497\
        );

    \I__2582\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11494\
        );

    \I__2581\ : Odrv12
    port map (
            O => \N__11497\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8EZ0\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__11494\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8EZ0\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__11489\,
            I => \N__11484\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__11488\,
            I => \N__11480\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__11487\,
            I => \N__11477\
        );

    \I__2576\ : InMux
    port map (
            O => \N__11484\,
            I => \N__11465\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11483\,
            I => \N__11465\
        );

    \I__2574\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11465\
        );

    \I__2573\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11465\
        );

    \I__2572\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11465\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__11465\,
            I => \Lab_UT.dspStr.cnt_fastZ0Z_2\
        );

    \I__2570\ : InMux
    port map (
            O => \N__11462\,
            I => \N__11459\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__11459\,
            I => \N__11452\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__11458\,
            I => \N__11449\
        );

    \I__2567\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11445\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11456\,
            I => \N__11440\
        );

    \I__2565\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11440\
        );

    \I__2564\ : Span4Mux_h
    port map (
            O => \N__11452\,
            I => \N__11437\
        );

    \I__2563\ : InMux
    port map (
            O => \N__11449\,
            I => \N__11432\
        );

    \I__2562\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11432\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__11445\,
            I => \N__11427\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__11440\,
            I => \N__11427\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__11437\,
            I => \Lab_UT_rx_data_0\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__11432\,
            I => \Lab_UT_rx_data_0\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__11427\,
            I => \Lab_UT_rx_data_0\
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__11420\,
            I => \N__11417\
        );

    \I__2555\ : InMux
    port map (
            O => \N__11417\,
            I => \N__11413\
        );

    \I__2554\ : InMux
    port map (
            O => \N__11416\,
            I => \N__11410\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__11413\,
            I => \N__11405\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__11410\,
            I => \N__11402\
        );

    \I__2551\ : InMux
    port map (
            O => \N__11409\,
            I => \N__11399\
        );

    \I__2550\ : InMux
    port map (
            O => \N__11408\,
            I => \N__11396\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__11405\,
            I => \Lab_UT_rx_data_1\
        );

    \I__2548\ : Odrv12
    port map (
            O => \N__11402\,
            I => \Lab_UT_rx_data_1\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__11399\,
            I => \Lab_UT_rx_data_1\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__11396\,
            I => \Lab_UT_rx_data_1\
        );

    \I__2545\ : InMux
    port map (
            O => \N__11387\,
            I => \N__11383\
        );

    \I__2544\ : InMux
    port map (
            O => \N__11386\,
            I => \N__11379\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__11383\,
            I => \N__11375\
        );

    \I__2542\ : InMux
    port map (
            O => \N__11382\,
            I => \N__11372\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__11379\,
            I => \N__11369\
        );

    \I__2540\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11366\
        );

    \I__2539\ : Odrv4
    port map (
            O => \N__11375\,
            I => \Lab_UT_rx_data_2\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__11372\,
            I => \Lab_UT_rx_data_2\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__11369\,
            I => \Lab_UT_rx_data_2\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__11366\,
            I => \Lab_UT_rx_data_2\
        );

    \I__2535\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11351\
        );

    \I__2534\ : InMux
    port map (
            O => \N__11356\,
            I => \N__11344\
        );

    \I__2533\ : InMux
    port map (
            O => \N__11355\,
            I => \N__11344\
        );

    \I__2532\ : InMux
    port map (
            O => \N__11354\,
            I => \N__11344\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__11351\,
            I => \N__11338\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__11344\,
            I => \N__11338\
        );

    \I__2529\ : InMux
    port map (
            O => \N__11343\,
            I => \N__11335\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__11338\,
            I => \Lab_UT_rx_data_3\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__11335\,
            I => \Lab_UT_rx_data_3\
        );

    \I__2526\ : InMux
    port map (
            O => \N__11330\,
            I => \N__11324\
        );

    \I__2525\ : InMux
    port map (
            O => \N__11329\,
            I => \N__11324\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__11324\,
            I => \N__11320\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__11323\,
            I => \N__11317\
        );

    \I__2522\ : Span4Mux_h
    port map (
            O => \N__11320\,
            I => \N__11314\
        );

    \I__2521\ : InMux
    port map (
            O => \N__11317\,
            I => \N__11311\
        );

    \I__2520\ : Odrv4
    port map (
            O => \N__11314\,
            I => \Lab_UT_rx_data_6\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__11311\,
            I => \Lab_UT_rx_data_6\
        );

    \I__2518\ : InMux
    port map (
            O => \N__11306\,
            I => \N__11303\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__11303\,
            I => \N__11300\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__11300\,
            I => \N__11295\
        );

    \I__2515\ : InMux
    port map (
            O => \N__11299\,
            I => \N__11290\
        );

    \I__2514\ : InMux
    port map (
            O => \N__11298\,
            I => \N__11290\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__11295\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9EZ0\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__11290\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9EZ0\
        );

    \I__2511\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11281\
        );

    \I__2510\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11273\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__11281\,
            I => \N__11270\
        );

    \I__2508\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11259\
        );

    \I__2507\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11259\
        );

    \I__2506\ : InMux
    port map (
            O => \N__11278\,
            I => \N__11259\
        );

    \I__2505\ : InMux
    port map (
            O => \N__11277\,
            I => \N__11259\
        );

    \I__2504\ : InMux
    port map (
            O => \N__11276\,
            I => \N__11259\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__11273\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__11270\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__11259\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__2500\ : InMux
    port map (
            O => \N__11252\,
            I => \N__11237\
        );

    \I__2499\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11237\
        );

    \I__2498\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11224\
        );

    \I__2497\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11224\
        );

    \I__2496\ : InMux
    port map (
            O => \N__11248\,
            I => \N__11224\
        );

    \I__2495\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11224\
        );

    \I__2494\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11224\
        );

    \I__2493\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11224\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__11244\,
            I => \N__11221\
        );

    \I__2491\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11214\
        );

    \I__2490\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11210\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__11237\,
            I => \N__11205\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__11224\,
            I => \N__11205\
        );

    \I__2487\ : InMux
    port map (
            O => \N__11221\,
            I => \N__11202\
        );

    \I__2486\ : InMux
    port map (
            O => \N__11220\,
            I => \N__11198\
        );

    \I__2485\ : InMux
    port map (
            O => \N__11219\,
            I => \N__11193\
        );

    \I__2484\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11193\
        );

    \I__2483\ : InMux
    port map (
            O => \N__11217\,
            I => \N__11190\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__11214\,
            I => \N__11187\
        );

    \I__2481\ : InMux
    port map (
            O => \N__11213\,
            I => \N__11184\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__11210\,
            I => \N__11180\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__11205\,
            I => \N__11175\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__11202\,
            I => \N__11175\
        );

    \I__2477\ : InMux
    port map (
            O => \N__11201\,
            I => \N__11172\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__11198\,
            I => \N__11169\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__11193\,
            I => \N__11166\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__11190\,
            I => \N__11161\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__11187\,
            I => \N__11161\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__11184\,
            I => \N__11158\
        );

    \I__2471\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11155\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__11180\,
            I => \N__11150\
        );

    \I__2469\ : Span4Mux_h
    port map (
            O => \N__11175\,
            I => \N__11150\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__11172\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__11169\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__2466\ : Odrv12
    port map (
            O => \N__11166\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__11161\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__11158\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__11155\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__11150\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__2460\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11129\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__11126\,
            I => \N__11123\
        );

    \I__2457\ : Span4Mux_h
    port map (
            O => \N__11123\,
            I => \N__11120\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__11120\,
            I => \uu2.mem0.w_addr_0\
        );

    \I__2455\ : CascadeMux
    port map (
            O => \N__11117\,
            I => \Lab_UT_L3_tx_data_0_5_cascade_\
        );

    \I__2454\ : InMux
    port map (
            O => \N__11114\,
            I => \N__11110\
        );

    \I__2453\ : InMux
    port map (
            O => \N__11113\,
            I => \N__11107\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__11110\,
            I => \Lab_UT_L3_tx_data_0_2_6\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__11107\,
            I => \Lab_UT_L3_tx_data_0_2_6\
        );

    \I__2450\ : InMux
    port map (
            O => \N__11102\,
            I => \N__11096\
        );

    \I__2449\ : InMux
    port map (
            O => \N__11101\,
            I => \N__11096\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__11096\,
            I => \N__11092\
        );

    \I__2447\ : InMux
    port map (
            O => \N__11095\,
            I => \N__11089\
        );

    \I__2446\ : Span4Mux_h
    port map (
            O => \N__11092\,
            I => \N__11083\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__11089\,
            I => \N__11080\
        );

    \I__2444\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11073\
        );

    \I__2443\ : InMux
    port map (
            O => \N__11087\,
            I => \N__11073\
        );

    \I__2442\ : InMux
    port map (
            O => \N__11086\,
            I => \N__11073\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__11083\,
            I => \uu2.un1_w_user_crZ0Z_4\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__11080\,
            I => \uu2.un1_w_user_crZ0Z_4\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__11073\,
            I => \uu2.un1_w_user_crZ0Z_4\
        );

    \I__2438\ : InMux
    port map (
            O => \N__11066\,
            I => \N__11063\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__11063\,
            I => \Lab_UT_L3_tx_data_0_2_1\
        );

    \I__2436\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11057\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__11057\,
            I => \Lab_UT_L3_tx_data_2_3\
        );

    \I__2434\ : InMux
    port map (
            O => \N__11054\,
            I => \N__11050\
        );

    \I__2433\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11047\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__11050\,
            I => \N__11043\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__11047\,
            I => \N__11040\
        );

    \I__2430\ : InMux
    port map (
            O => \N__11046\,
            I => \N__11037\
        );

    \I__2429\ : Odrv4
    port map (
            O => \N__11043\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87EZ0\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__11040\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87EZ0\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__11037\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87EZ0\
        );

    \I__2426\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11027\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__11027\,
            I => \N__11024\
        );

    \I__2424\ : Span4Mux_h
    port map (
            O => \N__11024\,
            I => \N__11020\
        );

    \I__2423\ : InMux
    port map (
            O => \N__11023\,
            I => \N__11017\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__11020\,
            I => \L3_tx_data_2\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__11017\,
            I => \L3_tx_data_2\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__11012\,
            I => \N__11009\
        );

    \I__2419\ : InMux
    port map (
            O => \N__11009\,
            I => \N__11002\
        );

    \I__2418\ : InMux
    port map (
            O => \N__11008\,
            I => \N__10993\
        );

    \I__2417\ : InMux
    port map (
            O => \N__11007\,
            I => \N__10993\
        );

    \I__2416\ : InMux
    port map (
            O => \N__11006\,
            I => \N__10993\
        );

    \I__2415\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10993\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__11002\,
            I => \Lab_UT.dspStr.cnt_fastZ0Z_1\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10993\,
            I => \Lab_UT.dspStr.cnt_fastZ0Z_1\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__10988\,
            I => \N__10981\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10970\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10970\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10970\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10984\,
            I => \N__10970\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10970\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10970\,
            I => \Lab_UT.dspStr.cnt_fastZ0Z_3\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10967\,
            I => \N__10964\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10964\,
            I => \N__10960\
        );

    \I__2403\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10957\
        );

    \I__2402\ : Odrv12
    port map (
            O => \N__10960\,
            I => \Lab_UT_L3_tx_data_0_4\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10957\,
            I => \Lab_UT_L3_tx_data_0_4\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10952\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_0\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10949\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_1\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10946\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_2\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10937\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10937\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10937\,
            I => \N__10932\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10936\,
            I => \N__10929\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10935\,
            I => \N__10926\
        );

    \I__2392\ : Span4Mux_v
    port map (
            O => \N__10932\,
            I => \N__10921\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10929\,
            I => \N__10911\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10926\,
            I => \N__10911\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10908\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10905\
        );

    \I__2387\ : Span4Mux_h
    port map (
            O => \N__10921\,
            I => \N__10902\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10895\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10895\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10918\,
            I => \N__10895\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10917\,
            I => \N__10890\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10890\
        );

    \I__2381\ : Span4Mux_h
    port map (
            O => \N__10911\,
            I => \N__10885\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__10908\,
            I => \N__10885\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10905\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__2378\ : Odrv4
    port map (
            O => \N__10902\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10895\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10890\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__10885\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10869\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__10873\,
            I => \N__10864\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__10872\,
            I => \N__10860\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10869\,
            I => \N__10856\
        );

    \I__2370\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10853\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10867\,
            I => \N__10850\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10864\,
            I => \N__10847\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10863\,
            I => \N__10840\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10840\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10840\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__10856\,
            I => \buart__rx_bitcount_3\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10853\,
            I => \buart__rx_bitcount_3\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10850\,
            I => \buart__rx_bitcount_3\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10847\,
            I => \buart__rx_bitcount_3\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__10840\,
            I => \buart__rx_bitcount_3\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__10829\,
            I => \N__10826\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10822\
        );

    \I__2357\ : InMux
    port map (
            O => \N__10825\,
            I => \N__10814\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10822\,
            I => \N__10811\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10821\,
            I => \N__10808\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10820\,
            I => \N__10799\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10819\,
            I => \N__10799\
        );

    \I__2352\ : InMux
    port map (
            O => \N__10818\,
            I => \N__10799\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10799\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10814\,
            I => \buart__rx_bitcount_2\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__10811\,
            I => \buart__rx_bitcount_2\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__10808\,
            I => \buart__rx_bitcount_2\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10799\,
            I => \buart__rx_bitcount_2\
        );

    \I__2346\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10787\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__2344\ : Span4Mux_v
    port map (
            O => \N__10784\,
            I => \N__10779\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10783\,
            I => \N__10774\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10782\,
            I => \N__10774\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__10779\,
            I => \N_87\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__10774\,
            I => \N_87\
        );

    \I__2339\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10766\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__10766\,
            I => \Lab_UT.rx_data_rdy\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10755\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10755\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10761\,
            I => \N__10749\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10760\,
            I => \N__10746\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__10755\,
            I => \N__10743\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10754\,
            I => \N__10740\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10753\,
            I => \N__10735\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10752\,
            I => \N__10735\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10749\,
            I => \buart__rx_bitcount_0\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10746\,
            I => \buart__rx_bitcount_0\
        );

    \I__2327\ : Odrv4
    port map (
            O => \N__10743\,
            I => \buart__rx_bitcount_0\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__10740\,
            I => \buart__rx_bitcount_0\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10735\,
            I => \buart__rx_bitcount_0\
        );

    \I__2324\ : InMux
    port map (
            O => \N__10724\,
            I => \N__10721\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10721\,
            I => \N__10718\
        );

    \I__2322\ : Span4Mux_h
    port map (
            O => \N__10718\,
            I => \N__10715\
        );

    \I__2321\ : Odrv4
    port map (
            O => \N__10715\,
            I => \resetGen.un3_reset_count_i_a3Z0Z_4\
        );

    \I__2320\ : InMux
    port map (
            O => \N__10712\,
            I => \N__10709\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__10709\,
            I => \N__10706\
        );

    \I__2318\ : Span4Mux_v
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__2317\ : Span4Mux_h
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__10700\,
            I => \Lab_UT_L3_tx_data_0_6\
        );

    \I__2315\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10692\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10686\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10695\,
            I => \N__10686\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__10692\,
            I => \N__10683\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__10691\,
            I => \N__10680\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__10686\,
            I => \N__10676\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__10683\,
            I => \N__10670\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10667\
        );

    \I__2307\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10661\
        );

    \I__2306\ : Span4Mux_v
    port map (
            O => \N__10676\,
            I => \N__10658\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10675\,
            I => \N__10655\
        );

    \I__2304\ : InMux
    port map (
            O => \N__10674\,
            I => \N__10650\
        );

    \I__2303\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10650\
        );

    \I__2302\ : Span4Mux_h
    port map (
            O => \N__10670\,
            I => \N__10645\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10667\,
            I => \N__10645\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10638\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10638\
        );

    \I__2298\ : InMux
    port map (
            O => \N__10664\,
            I => \N__10638\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__10661\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__10658\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__10655\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__10650\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__2293\ : Odrv4
    port map (
            O => \N__10645\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__10638\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__10625\,
            I => \N__10621\
        );

    \I__2290\ : CascadeMux
    port map (
            O => \N__10624\,
            I => \N__10614\
        );

    \I__2289\ : InMux
    port map (
            O => \N__10621\,
            I => \N__10610\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__10620\,
            I => \N__10607\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__10619\,
            I => \N__10604\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__10618\,
            I => \N__10601\
        );

    \I__2285\ : InMux
    port map (
            O => \N__10617\,
            I => \N__10596\
        );

    \I__2284\ : InMux
    port map (
            O => \N__10614\,
            I => \N__10596\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__10613\,
            I => \N__10592\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__10610\,
            I => \N__10588\
        );

    \I__2281\ : InMux
    port map (
            O => \N__10607\,
            I => \N__10583\
        );

    \I__2280\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10583\
        );

    \I__2279\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10580\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__10596\,
            I => \N__10575\
        );

    \I__2277\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10568\
        );

    \I__2276\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10568\
        );

    \I__2275\ : InMux
    port map (
            O => \N__10591\,
            I => \N__10568\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__10588\,
            I => \N__10563\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__10583\,
            I => \N__10563\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__10580\,
            I => \N__10560\
        );

    \I__2271\ : InMux
    port map (
            O => \N__10579\,
            I => \N__10557\
        );

    \I__2270\ : InMux
    port map (
            O => \N__10578\,
            I => \N__10554\
        );

    \I__2269\ : Span4Mux_v
    port map (
            O => \N__10575\,
            I => \N__10549\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__10568\,
            I => \N__10549\
        );

    \I__2267\ : Span4Mux_h
    port map (
            O => \N__10563\,
            I => \N__10546\
        );

    \I__2266\ : Span4Mux_h
    port map (
            O => \N__10560\,
            I => \N__10543\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__10557\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10554\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__10549\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__10546\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__10543\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__2260\ : InMux
    port map (
            O => \N__10532\,
            I => \N__10529\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__10529\,
            I => \buart.Z_tx.bitcount_RNO_0Z0Z_2\
        );

    \I__2258\ : InMux
    port map (
            O => \N__10526\,
            I => \buart.Z_tx.un1_bitcount_cry_1\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__10523\,
            I => \N__10520\
        );

    \I__2256\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10513\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__10519\,
            I => \N__10510\
        );

    \I__2254\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10500\
        );

    \I__2253\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10500\
        );

    \I__2252\ : InMux
    port map (
            O => \N__10516\,
            I => \N__10497\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__10513\,
            I => \N__10494\
        );

    \I__2250\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10489\
        );

    \I__2249\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10489\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__10508\,
            I => \N__10481\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__10507\,
            I => \N__10478\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__10506\,
            I => \N__10473\
        );

    \I__2245\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10466\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__10500\,
            I => \N__10457\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__10497\,
            I => \N__10457\
        );

    \I__2242\ : Span4Mux_h
    port map (
            O => \N__10494\,
            I => \N__10457\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__10489\,
            I => \N__10457\
        );

    \I__2240\ : InMux
    port map (
            O => \N__10488\,
            I => \N__10450\
        );

    \I__2239\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10450\
        );

    \I__2238\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10450\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10485\,
            I => \N__10445\
        );

    \I__2236\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10445\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10438\
        );

    \I__2234\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10438\
        );

    \I__2233\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10438\
        );

    \I__2232\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10431\
        );

    \I__2231\ : InMux
    port map (
            O => \N__10473\,
            I => \N__10431\
        );

    \I__2230\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10431\
        );

    \I__2229\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10424\
        );

    \I__2228\ : InMux
    port map (
            O => \N__10470\,
            I => \N__10424\
        );

    \I__2227\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10424\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__10466\,
            I => \N__10421\
        );

    \I__2225\ : Span4Mux_h
    port map (
            O => \N__10457\,
            I => \N__10418\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__10450\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__10445\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__10438\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__10431\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__10424\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2219\ : Odrv12
    port map (
            O => \N__10421\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__10418\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2217\ : InMux
    port map (
            O => \N__10403\,
            I => \buart.Z_tx.un1_bitcount_cry_2\
        );

    \I__2216\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__10397\,
            I => \buart.Z_tx.bitcount_RNIM5O32Z0Z_2\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__10394\,
            I => \N__10390\
        );

    \I__2213\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10384\
        );

    \I__2212\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10384\
        );

    \I__2211\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10381\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__10384\,
            I => \N__10376\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__10381\,
            I => \N__10376\
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__10376\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__10373\,
            I => \N__10368\
        );

    \I__2206\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10362\
        );

    \I__2205\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10362\
        );

    \I__2204\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10357\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10357\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__10362\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__10357\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__2199\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10344\
        );

    \I__2198\ : InMux
    port map (
            O => \N__10348\,
            I => \N__10339\
        );

    \I__2197\ : InMux
    port map (
            O => \N__10347\,
            I => \N__10339\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__10344\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__10339\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__10334\,
            I => \buart__tx_uart_busy_0_cascade_\
        );

    \I__2193\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__10328\,
            I => \buart.Z_tx.bitcount_RNIL4O32Z0Z_1\
        );

    \I__2191\ : InMux
    port map (
            O => \N__10325\,
            I => \N__10310\
        );

    \I__2190\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10310\
        );

    \I__2189\ : InMux
    port map (
            O => \N__10323\,
            I => \N__10310\
        );

    \I__2188\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10303\
        );

    \I__2187\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10303\
        );

    \I__2186\ : InMux
    port map (
            O => \N__10320\,
            I => \N__10303\
        );

    \I__2185\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10296\
        );

    \I__2184\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10296\
        );

    \I__2183\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10296\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__10310\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__10303\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__10296\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__10289\,
            I => \N__10281\
        );

    \I__2178\ : InMux
    port map (
            O => \N__10288\,
            I => \N__10265\
        );

    \I__2177\ : InMux
    port map (
            O => \N__10287\,
            I => \N__10265\
        );

    \I__2176\ : InMux
    port map (
            O => \N__10286\,
            I => \N__10265\
        );

    \I__2175\ : InMux
    port map (
            O => \N__10285\,
            I => \N__10265\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__10284\,
            I => \N__10262\
        );

    \I__2173\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10259\
        );

    \I__2172\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10254\
        );

    \I__2171\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10254\
        );

    \I__2170\ : InMux
    port map (
            O => \N__10278\,
            I => \N__10245\
        );

    \I__2169\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10245\
        );

    \I__2168\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10245\
        );

    \I__2167\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10245\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__10274\,
            I => \N__10241\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__10265\,
            I => \N__10233\
        );

    \I__2164\ : InMux
    port map (
            O => \N__10262\,
            I => \N__10230\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__10259\,
            I => \N__10223\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__10254\,
            I => \N__10223\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__10245\,
            I => \N__10223\
        );

    \I__2160\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10216\
        );

    \I__2159\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10216\
        );

    \I__2158\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10216\
        );

    \I__2157\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10207\
        );

    \I__2156\ : InMux
    port map (
            O => \N__10238\,
            I => \N__10207\
        );

    \I__2155\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10207\
        );

    \I__2154\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10207\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__10233\,
            I => \N__10204\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__10230\,
            I => \buart__tx_uart_busy_0\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__10223\,
            I => \buart__tx_uart_busy_0\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__10216\,
            I => \buart__tx_uart_busy_0\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__10207\,
            I => \buart__tx_uart_busy_0\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__10204\,
            I => \buart__tx_uart_busy_0\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__10193\,
            I => \N__10189\
        );

    \I__2146\ : InMux
    port map (
            O => \N__10192\,
            I => \N__10186\
        );

    \I__2145\ : InMux
    port map (
            O => \N__10189\,
            I => \N__10183\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__10186\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__10183\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__2142\ : InMux
    port map (
            O => \N__10178\,
            I => \N__10175\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__10175\,
            I => \buart.Z_tx.un1_bitcount_axb_3\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__10172\,
            I => \N__10169\
        );

    \I__2139\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10165\
        );

    \I__2138\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10162\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__10165\,
            I => \N__10159\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__10162\,
            I => \Lab_UT.dspStr.cnt11_0_i\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__10159\,
            I => \Lab_UT.dspStr.cnt11_0_i\
        );

    \I__2134\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10151\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__10151\,
            I => \N__10148\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__10148\,
            I => \N__10145\
        );

    \I__2131\ : Span4Mux_h
    port map (
            O => \N__10145\,
            I => \N__10140\
        );

    \I__2130\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10137\
        );

    \I__2129\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10134\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__10140\,
            I => \Lab_UT.dspStr.cntZ0Z_0\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__10137\,
            I => \Lab_UT.dspStr.cntZ0Z_0\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__10134\,
            I => \Lab_UT.dspStr.cntZ0Z_0\
        );

    \I__2125\ : InMux
    port map (
            O => \N__10127\,
            I => \Lab_UT.didpuu0.didpsones.un1_q_cry_0\
        );

    \I__2124\ : InMux
    port map (
            O => \N__10124\,
            I => \N__10121\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__10121\,
            I => \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_2\
        );

    \I__2122\ : InMux
    port map (
            O => \N__10118\,
            I => \Lab_UT.didpuu0.didpsones.un1_q_cry_1\
        );

    \I__2121\ : InMux
    port map (
            O => \N__10115\,
            I => \Lab_UT.didpuu0.didpsones.un1_q_cry_2\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__10112\,
            I => \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_3_cascade_\
        );

    \I__2119\ : InMux
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__10106\,
            I => \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_0\
        );

    \I__2117\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10100\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__10100\,
            I => \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_1\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__10097\,
            I => \N__10092\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__10096\,
            I => \N__10089\
        );

    \I__2113\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10082\
        );

    \I__2112\ : InMux
    port map (
            O => \N__10092\,
            I => \N__10082\
        );

    \I__2111\ : InMux
    port map (
            O => \N__10089\,
            I => \N__10082\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__10082\,
            I => \Lab_UT.didpuu0.didpsones.q13_0\
        );

    \I__2109\ : InMux
    port map (
            O => \N__10079\,
            I => \N__10069\
        );

    \I__2108\ : InMux
    port map (
            O => \N__10078\,
            I => \N__10069\
        );

    \I__2107\ : InMux
    port map (
            O => \N__10077\,
            I => \N__10069\
        );

    \I__2106\ : InMux
    port map (
            O => \N__10076\,
            I => \N__10066\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__10069\,
            I => \N__10060\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__10066\,
            I => \N__10060\
        );

    \I__2103\ : InMux
    port map (
            O => \N__10065\,
            I => \N__10056\
        );

    \I__2102\ : Span4Mux_h
    port map (
            O => \N__10060\,
            I => \N__10053\
        );

    \I__2101\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10050\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__10056\,
            I => \N__10047\
        );

    \I__2099\ : Span4Mux_v
    port map (
            O => \N__10053\,
            I => \N__10044\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__10050\,
            I => \N__10039\
        );

    \I__2097\ : Span4Mux_h
    port map (
            O => \N__10047\,
            I => \N__10039\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__10044\,
            I => rst
        );

    \I__2095\ : Odrv4
    port map (
            O => \N__10039\,
            I => rst
        );

    \I__2094\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10031\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__10031\,
            I => \buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0\
        );

    \I__2092\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10025\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__10025\,
            I => \buart.Z_tx.bitcount_RNO_0Z0Z_1\
        );

    \I__2090\ : InMux
    port map (
            O => \N__10022\,
            I => \buart.Z_tx.un1_bitcount_cry_0\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__10019\,
            I => \N__10015\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__10018\,
            I => \N__10011\
        );

    \I__2087\ : InMux
    port map (
            O => \N__10015\,
            I => \N__10008\
        );

    \I__2086\ : InMux
    port map (
            O => \N__10014\,
            I => \N__10002\
        );

    \I__2085\ : InMux
    port map (
            O => \N__10011\,
            I => \N__9999\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__10008\,
            I => \N__9996\
        );

    \I__2083\ : InMux
    port map (
            O => \N__10007\,
            I => \N__9989\
        );

    \I__2082\ : InMux
    port map (
            O => \N__10006\,
            I => \N__9989\
        );

    \I__2081\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9989\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__10002\,
            I => \uu2.w_addr_displaying_fastZ0Z_4\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9999\,
            I => \uu2.w_addr_displaying_fastZ0Z_4\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__9996\,
            I => \uu2.w_addr_displaying_fastZ0Z_4\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__9989\,
            I => \uu2.w_addr_displaying_fastZ0Z_4\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9977\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__9974\,
            I => \uu2.mem0.Z_decfrac105_7_3_2\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__9971\,
            I => \uu2.w_addr_displaying_4_8_cascade_\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__9968\,
            I => \N__9961\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9958\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__9966\,
            I => \N__9954\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9951\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9946\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9946\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9958\,
            I => \N__9940\
        );

    \I__2065\ : InMux
    port map (
            O => \N__9957\,
            I => \N__9937\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9954\,
            I => \N__9934\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__9951\,
            I => \N__9929\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9946\,
            I => \N__9929\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9922\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9922\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9943\,
            I => \N__9922\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__9940\,
            I => \N__9917\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__9937\,
            I => \N__9917\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__9934\,
            I => \N__9914\
        );

    \I__2055\ : Span4Mux_v
    port map (
            O => \N__9929\,
            I => \N__9911\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__9922\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__9917\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__9914\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__9911\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9896\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9893\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9900\,
            I => \N__9888\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9899\,
            I => \N__9888\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__9896\,
            I => \N__9885\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__9893\,
            I => \N__9880\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9888\,
            I => \N__9880\
        );

    \I__2043\ : Odrv12
    port map (
            O => \N__9885\,
            I => \uu2.un15_w_data_displaying\
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__9880\,
            I => \uu2.un15_w_data_displaying\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__9875\,
            I => \uu2.un15_w_data_displaying_cascade_\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__9872\,
            I => \N__9866\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__9871\,
            I => \N__9862\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9858\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9855\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9866\,
            I => \N__9852\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9865\,
            I => \N__9849\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9862\,
            I => \N__9844\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9861\,
            I => \N__9844\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9858\,
            I => \N__9839\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9855\,
            I => \N__9834\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__9852\,
            I => \N__9834\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9849\,
            I => \N__9829\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9844\,
            I => \N__9829\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9826\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9823\
        );

    \I__2025\ : Span4Mux_v
    port map (
            O => \N__9839\,
            I => \N__9820\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__9834\,
            I => \N__9817\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__9829\,
            I => \N__9814\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__9826\,
            I => \N__9811\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9823\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__9820\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__9817\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__9814\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__9811\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9800\,
            I => \N__9797\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9797\,
            I => \N__9792\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9789\
        );

    \I__2013\ : InMux
    port map (
            O => \N__9795\,
            I => \N__9784\
        );

    \I__2012\ : Span4Mux_h
    port map (
            O => \N__9792\,
            I => \N__9781\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9789\,
            I => \N__9778\
        );

    \I__2010\ : InMux
    port map (
            O => \N__9788\,
            I => \N__9773\
        );

    \I__2009\ : InMux
    port map (
            O => \N__9787\,
            I => \N__9773\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9784\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__9781\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__2006\ : Odrv4
    port map (
            O => \N__9778\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9773\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__9764\,
            I => \N__9757\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__9763\,
            I => \N__9754\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__9762\,
            I => \N__9751\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__9761\,
            I => \N__9746\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__9760\,
            I => \N__9743\
        );

    \I__1999\ : InMux
    port map (
            O => \N__9757\,
            I => \N__9738\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9738\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9751\,
            I => \N__9731\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9750\,
            I => \N__9731\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9731\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9746\,
            I => \N__9726\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9726\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__9738\,
            I => \N__9723\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__9731\,
            I => \N__9718\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__9726\,
            I => \N__9718\
        );

    \I__1989\ : Span4Mux_v
    port map (
            O => \N__9723\,
            I => \N__9715\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__9718\,
            I => \N__9712\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__9715\,
            I => \uu2.un448_ci_5\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__9712\,
            I => \uu2.un448_ci_5\
        );

    \I__1985\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9700\
        );

    \I__1984\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9696\
        );

    \I__1983\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9692\
        );

    \I__1982\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9689\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__9703\,
            I => \N__9685\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__9700\,
            I => \N__9682\
        );

    \I__1979\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9679\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__9696\,
            I => \N__9676\
        );

    \I__1977\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9673\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__9692\,
            I => \N__9664\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__9689\,
            I => \N__9664\
        );

    \I__1974\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9659\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9685\,
            I => \N__9659\
        );

    \I__1972\ : Span4Mux_v
    port map (
            O => \N__9682\,
            I => \N__9654\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__9679\,
            I => \N__9654\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__9676\,
            I => \N__9649\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__9673\,
            I => \N__9649\
        );

    \I__1968\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9640\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9671\,
            I => \N__9640\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9640\
        );

    \I__1965\ : InMux
    port map (
            O => \N__9669\,
            I => \N__9640\
        );

    \I__1964\ : Span4Mux_v
    port map (
            O => \N__9664\,
            I => \N__9637\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__9659\,
            I => \N__9634\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__9654\,
            I => \N__9631\
        );

    \I__1961\ : Span4Mux_v
    port map (
            O => \N__9649\,
            I => \N__9628\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__9640\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__9637\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__9634\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__9631\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__9628\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__1955\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9608\
        );

    \I__1954\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9608\
        );

    \I__1953\ : InMux
    port map (
            O => \N__9615\,
            I => \N__9608\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__9608\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9599\
        );

    \I__1950\ : InMux
    port map (
            O => \N__9604\,
            I => \N__9590\
        );

    \I__1949\ : InMux
    port map (
            O => \N__9603\,
            I => \N__9590\
        );

    \I__1948\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9590\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__9599\,
            I => \N__9586\
        );

    \I__1946\ : InMux
    port map (
            O => \N__9598\,
            I => \N__9583\
        );

    \I__1945\ : InMux
    port map (
            O => \N__9597\,
            I => \N__9578\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__9590\,
            I => \N__9575\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9572\
        );

    \I__1942\ : Span4Mux_v
    port map (
            O => \N__9586\,
            I => \N__9567\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__9583\,
            I => \N__9567\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9582\,
            I => \N__9564\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9561\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__9578\,
            I => \N__9556\
        );

    \I__1937\ : Span4Mux_h
    port map (
            O => \N__9575\,
            I => \N__9556\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__9572\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__9567\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__9564\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__9561\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__9556\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__1931\ : InMux
    port map (
            O => \N__9545\,
            I => \N__9541\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__9544\,
            I => \N__9535\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__9541\,
            I => \N__9531\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9528\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__9539\,
            I => \N__9524\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9538\,
            I => \N__9519\
        );

    \I__1925\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9516\
        );

    \I__1924\ : InMux
    port map (
            O => \N__9534\,
            I => \N__9513\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__9531\,
            I => \N__9510\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9528\,
            I => \N__9507\
        );

    \I__1921\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9504\
        );

    \I__1920\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9497\
        );

    \I__1919\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9497\
        );

    \I__1918\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9497\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__9519\,
            I => \N__9494\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__9516\,
            I => \N__9489\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__9513\,
            I => \N__9489\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__9510\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__9507\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__9504\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__9497\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__9494\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__9489\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__1908\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9473\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__9473\,
            I => \uu2.mem0.bitmap_pmux_1_1_i_a5_1_0\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__9470\,
            I => \uu2.mem0.g1_1_0_cascade_\
        );

    \I__1905\ : InMux
    port map (
            O => \N__9467\,
            I => \N__9464\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__9464\,
            I => \N__9459\
        );

    \I__1903\ : InMux
    port map (
            O => \N__9463\,
            I => \N__9456\
        );

    \I__1902\ : InMux
    port map (
            O => \N__9462\,
            I => \N__9453\
        );

    \I__1901\ : Span4Mux_h
    port map (
            O => \N__9459\,
            I => \N__9448\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__9456\,
            I => \N__9448\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__9453\,
            I => \N__9445\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__9448\,
            I => \uu2.Z_decfrac106_5\
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__9445\,
            I => \uu2.Z_decfrac106_5\
        );

    \I__1896\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__1894\ : Span12Mux_s7_h
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__1893\ : Odrv12
    port map (
            O => \N__9431\,
            I => \uu2.mem0.g0_2_0\
        );

    \I__1892\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9425\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__9425\,
            I => \uu2.mem0.bitmap_pmux_1_1_i_a5_2_3_1_0\
        );

    \I__1890\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9416\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__9421\,
            I => \N__9413\
        );

    \I__1888\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9406\
        );

    \I__1887\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9403\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__9416\,
            I => \N__9400\
        );

    \I__1885\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9397\
        );

    \I__1884\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9392\
        );

    \I__1883\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9392\
        );

    \I__1882\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9389\
        );

    \I__1881\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9386\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__9406\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__9403\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__9400\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__9397\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__9392\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__9389\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__9386\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1873\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9362\
        );

    \I__1872\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9362\
        );

    \I__1871\ : InMux
    port map (
            O => \N__9369\,
            I => \N__9362\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__9362\,
            I => \N__9358\
        );

    \I__1869\ : InMux
    port map (
            O => \N__9361\,
            I => \N__9355\
        );

    \I__1868\ : Span4Mux_h
    port map (
            O => \N__9358\,
            I => \N__9352\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__9355\,
            I => \N__9349\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__9352\,
            I => \uu2.Z_decfrac105_7_2\
        );

    \I__1865\ : Odrv4
    port map (
            O => \N__9349\,
            I => \uu2.Z_decfrac105_7_2\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__9344\,
            I => \N__9339\
        );

    \I__1863\ : InMux
    port map (
            O => \N__9343\,
            I => \N__9331\
        );

    \I__1862\ : InMux
    port map (
            O => \N__9342\,
            I => \N__9331\
        );

    \I__1861\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9331\
        );

    \I__1860\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9328\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__9331\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__9328\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__9323\,
            I => \L3_tx_data_0_cascade_\
        );

    \I__1856\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9317\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__9317\,
            I => \N__9314\
        );

    \I__1854\ : Span4Mux_h
    port map (
            O => \N__9314\,
            I => \N__9308\
        );

    \I__1853\ : InMux
    port map (
            O => \N__9313\,
            I => \N__9301\
        );

    \I__1852\ : InMux
    port map (
            O => \N__9312\,
            I => \N__9301\
        );

    \I__1851\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9301\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__9308\,
            I => \uu2.un1_w_user_crZ0Z_1\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__9301\,
            I => \uu2.un1_w_user_crZ0Z_1\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__9296\,
            I => \uu2.w_addr_displaying_RNIQKOV8Z0Z_8_cascade_\
        );

    \I__1847\ : InMux
    port map (
            O => \N__9293\,
            I => \N__9281\
        );

    \I__1846\ : InMux
    port map (
            O => \N__9292\,
            I => \N__9281\
        );

    \I__1845\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9281\
        );

    \I__1844\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9281\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__9281\,
            I => \N__9276\
        );

    \I__1842\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9273\
        );

    \I__1841\ : InMux
    port map (
            O => \N__9279\,
            I => \N__9270\
        );

    \I__1840\ : Span4Mux_h
    port map (
            O => \N__9276\,
            I => \N__9267\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__9273\,
            I => \L3_tx_data_rdy\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__9270\,
            I => \L3_tx_data_rdy\
        );

    \I__1837\ : Odrv4
    port map (
            O => \N__9267\,
            I => \L3_tx_data_rdy\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__9260\,
            I => \uu2.un21_w_addr_displaying_i_cascade_\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__1834\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__1832\ : Span4Mux_h
    port map (
            O => \N__9248\,
            I => \N__9245\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__9245\,
            I => \uu2.mem0.g0_i_a11_1_0\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__9242\,
            I => \N__9239\
        );

    \I__1829\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9232\
        );

    \I__1828\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9229\
        );

    \I__1827\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9225\
        );

    \I__1826\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9220\
        );

    \I__1825\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9220\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__9232\,
            I => \N__9217\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__9229\,
            I => \N__9214\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__9228\,
            I => \N__9211\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__9225\,
            I => \N__9206\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__9220\,
            I => \N__9199\
        );

    \I__1819\ : Span4Mux_h
    port map (
            O => \N__9217\,
            I => \N__9199\
        );

    \I__1818\ : Span4Mux_h
    port map (
            O => \N__9214\,
            I => \N__9196\
        );

    \I__1817\ : InMux
    port map (
            O => \N__9211\,
            I => \N__9193\
        );

    \I__1816\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9188\
        );

    \I__1815\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9188\
        );

    \I__1814\ : Span4Mux_v
    port map (
            O => \N__9206\,
            I => \N__9185\
        );

    \I__1813\ : InMux
    port map (
            O => \N__9205\,
            I => \N__9180\
        );

    \I__1812\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9180\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__9199\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__9196\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__9193\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__9188\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__9185\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__9180\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__9167\,
            I => \uu2.mem0.g3_0_cascade_\
        );

    \I__1804\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9157\
        );

    \I__1803\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9157\
        );

    \I__1802\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9152\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__9157\,
            I => \N__9149\
        );

    \I__1800\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9145\
        );

    \I__1799\ : InMux
    port map (
            O => \N__9155\,
            I => \N__9142\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__9152\,
            I => \N__9139\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__9149\,
            I => \N__9129\
        );

    \I__1796\ : InMux
    port map (
            O => \N__9148\,
            I => \N__9126\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__9145\,
            I => \N__9123\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__9142\,
            I => \N__9120\
        );

    \I__1793\ : Span4Mux_h
    port map (
            O => \N__9139\,
            I => \N__9117\
        );

    \I__1792\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9110\
        );

    \I__1791\ : InMux
    port map (
            O => \N__9137\,
            I => \N__9110\
        );

    \I__1790\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9110\
        );

    \I__1789\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9103\
        );

    \I__1788\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9103\
        );

    \I__1787\ : InMux
    port map (
            O => \N__9133\,
            I => \N__9103\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9132\,
            I => \N__9100\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__9129\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__9126\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1783\ : Odrv4
    port map (
            O => \N__9123\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__9120\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__9117\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__9110\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__9103\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__9100\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1777\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__1775\ : Odrv4
    port map (
            O => \N__9077\,
            I => \uu2.mem0.un1_segment4_0_i_i_0_0\
        );

    \I__1774\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9071\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__9071\,
            I => \N__9068\
        );

    \I__1772\ : Odrv12
    port map (
            O => \N__9068\,
            I => \uu2.mem0.g0_i_a11_3_1\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__9065\,
            I => \uu2.mem0.g0_i_a11_7_1_cascade_\
        );

    \I__1770\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__9056\,
            I => \uu2.mem0.g0_i_5_1\
        );

    \I__1767\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9047\
        );

    \I__1766\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9040\
        );

    \I__1765\ : InMux
    port map (
            O => \N__9051\,
            I => \N__9040\
        );

    \I__1764\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9040\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__9047\,
            I => \Lab_UT_dspStr_cnt_1_rep1\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__9040\,
            I => \Lab_UT_dspStr_cnt_1_rep1\
        );

    \I__1761\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__9032\,
            I => \N__9029\
        );

    \I__1759\ : Span4Mux_h
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__1758\ : Odrv4
    port map (
            O => \N__9026\,
            I => \Lab_UT_dspStr_un36_dOut\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__9023\,
            I => \Lab_UT_dspStr_un36_dOut_cascade_\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__9020\,
            I => \uu2.un27_N_6_mux_cascade_\
        );

    \I__1755\ : InMux
    port map (
            O => \N__9017\,
            I => \N__9014\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__9014\,
            I => \N__9011\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__9011\,
            I => \uu2.un27_w_addr_user_iZ0Z_1\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__9008\,
            I => \N__9003\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__9007\,
            I => \N__9000\
        );

    \I__1750\ : InMux
    port map (
            O => \N__9006\,
            I => \N__8996\
        );

    \I__1749\ : InMux
    port map (
            O => \N__9003\,
            I => \N__8989\
        );

    \I__1748\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8989\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8989\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8996\,
            I => \Lab_UT_dspStr_cnt_3_rep1\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8989\,
            I => \Lab_UT_dspStr_cnt_3_rep1\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8975\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8983\,
            I => \N__8975\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8982\,
            I => \N__8968\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8968\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8968\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8975\,
            I => \Lab_UT_dspStr_cnt_2_rep1\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__8968\,
            I => \Lab_UT_dspStr_cnt_2_rep1\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8960\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__8960\,
            I => \N__8956\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__8959\,
            I => \N__8953\
        );

    \I__1734\ : Span4Mux_h
    port map (
            O => \N__8956\,
            I => \N__8950\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8953\,
            I => \N__8947\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__8950\,
            I => \L3_tx_data_0\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__8947\,
            I => \L3_tx_data_0\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8939\,
            I => \uu2.w_m5_i_a3Z0Z_2\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8933\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8933\,
            I => \Lab_UT.dictrluu0.dek.det_NZ0Z_4\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__8930\,
            I => \uu2.un1_w_user_lf_0_0Z0Z_0_cascade_\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8924\,
            I => \uu2.un1_w_user_lf_2\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__8918\,
            I => \N__8914\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8917\,
            I => \N__8911\
        );

    \I__1720\ : Span4Mux_v
    port map (
            O => \N__8914\,
            I => \N__8908\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8911\,
            I => \uu2.un2_w_addr_user\
        );

    \I__1718\ : Odrv4
    port map (
            O => \N__8908\,
            I => \uu2.un2_w_addr_user\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__8903\,
            I => \uu2.un1_w_user_lf_2_cascade_\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8897\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8897\,
            I => \uu2.un27_N_6_mux_0\
        );

    \I__1714\ : IoInMux
    port map (
            O => \N__8894\,
            I => \N__8889\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8886\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__8892\,
            I => \N__8883\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8889\,
            I => \N__8880\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8886\,
            I => \N__8877\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8874\
        );

    \I__1708\ : Span4Mux_s2_v
    port map (
            O => \N__8880\,
            I => \N__8871\
        );

    \I__1707\ : Span4Mux_h
    port map (
            O => \N__8877\,
            I => \N__8866\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8874\,
            I => \N__8866\
        );

    \I__1705\ : Span4Mux_h
    port map (
            O => \N__8871\,
            I => \N__8863\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__8866\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__8863\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__8858\,
            I => \uu2.w_addr_user_RNILDNK6Z0Z_4_cascade_\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8848\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8848\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8839\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8848\,
            I => \N__8836\
        );

    \I__1697\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8829\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8829\
        );

    \I__1695\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8829\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8822\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8822\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8822\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__8839\,
            I => \N__8819\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__8836\,
            I => \uu2.un27_w_addr_user_i\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8829\,
            I => \uu2.un27_w_addr_user_i\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8822\,
            I => \uu2.un27_w_addr_user_i\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__8819\,
            I => \uu2.un27_w_addr_user_i\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__8810\,
            I => \uu2.un1_w_user_lf_5_a0Z0Z_5_cascade_\
        );

    \I__1685\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8804\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__8804\,
            I => \N__8800\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8797\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__8800\,
            I => \uu2.un1_w_user_lf_5_aZ0Z0\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__8797\,
            I => \uu2.un1_w_user_lf_5_aZ0Z0\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__8792\,
            I => \uu2.w_addr_user_2Z0Z_1_cascade_\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__8789\,
            I => \uu2.w_addr_userZ2Z_1_cascade_\
        );

    \I__1678\ : SRMux
    port map (
            O => \N__8786\,
            I => \N__8782\
        );

    \I__1677\ : SRMux
    port map (
            O => \N__8785\,
            I => \N__8778\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__8782\,
            I => \N__8774\
        );

    \I__1675\ : SRMux
    port map (
            O => \N__8781\,
            I => \N__8771\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8778\,
            I => \N__8768\
        );

    \I__1673\ : SRMux
    port map (
            O => \N__8777\,
            I => \N__8765\
        );

    \I__1672\ : Span4Mux_h
    port map (
            O => \N__8774\,
            I => \N__8762\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__8771\,
            I => \N__8755\
        );

    \I__1670\ : Span4Mux_s3_v
    port map (
            O => \N__8768\,
            I => \N__8755\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8765\,
            I => \N__8755\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__8762\,
            I => \uu2.w_addr_user_RNIT1MGDZ0Z_4\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__8755\,
            I => \uu2.w_addr_user_RNIT1MGDZ0Z_4\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8747\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8747\,
            I => \uu2.w_addr_user_1_0\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__8744\,
            I => \Lab_UT.dictrluu0.dek.det_NZ0Z_5_cascade_\
        );

    \I__1663\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8738\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__8735\,
            I => \N__8732\
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__8732\,
            I => \uu2.mem0.N_1476_0_0_0\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__8726\,
            I => \Lab_UT.dspStr.cnt11_1\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8723\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8720\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__1655\ : InMux
    port map (
            O => \N__8717\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__1654\ : InMux
    port map (
            O => \N__8714\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__1653\ : InMux
    port map (
            O => \N__8711\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__8708\,
            I => \N__8705\
        );

    \I__1651\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8699\
        );

    \I__1650\ : InMux
    port map (
            O => \N__8704\,
            I => \N__8699\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__8699\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8687\
        );

    \I__1646\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8687\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__8687\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__8684\,
            I => \N__8680\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8683\,
            I => \N__8677\
        );

    \I__1642\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8674\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8677\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__8674\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__1639\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8663\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8668\,
            I => \N__8663\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__8663\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__8660\,
            I => \N__8656\
        );

    \I__1635\ : InMux
    port map (
            O => \N__8659\,
            I => \N__8652\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8649\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8646\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__8652\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__8649\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__8646\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8631\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8638\,
            I => \N__8631\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8637\,
            I => \N__8628\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8636\,
            I => \N__8625\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8631\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__8628\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8625\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__8618\,
            I => \N__8614\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__8617\,
            I => \N__8611\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8606\
        );

    \I__1619\ : InMux
    port map (
            O => \N__8611\,
            I => \N__8606\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__8606\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8603\,
            I => \N__8600\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__8600\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__8597\,
            I => \Lab_UT.didpuu0.didpsones.q13_0_cascade_\
        );

    \I__1614\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__8591\,
            I => \uu2.g0_3Z0Z_0\
        );

    \I__1612\ : CEMux
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8585\,
            I => \N__8580\
        );

    \I__1610\ : CEMux
    port map (
            O => \N__8584\,
            I => \N__8577\
        );

    \I__1609\ : CEMux
    port map (
            O => \N__8583\,
            I => \N__8574\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__8580\,
            I => \N__8571\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__8577\,
            I => \N__8568\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__8574\,
            I => \N__8565\
        );

    \I__1605\ : Span4Mux_h
    port map (
            O => \N__8571\,
            I => \N__8562\
        );

    \I__1604\ : Span4Mux_h
    port map (
            O => \N__8568\,
            I => \N__8559\
        );

    \I__1603\ : Span4Mux_h
    port map (
            O => \N__8565\,
            I => \N__8556\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__8562\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__8559\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__8556\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8543\
        );

    \I__1598\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8538\
        );

    \I__1597\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8538\
        );

    \I__1596\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8535\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8543\,
            I => \N__8529\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__8538\,
            I => \N__8529\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__8535\,
            I => \N__8526\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__8534\,
            I => \N__8522\
        );

    \I__1591\ : Span4Mux_h
    port map (
            O => \N__8529\,
            I => \N__8517\
        );

    \I__1590\ : Span4Mux_h
    port map (
            O => \N__8526\,
            I => \N__8514\
        );

    \I__1589\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8511\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8506\
        );

    \I__1587\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8506\
        );

    \I__1586\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8503\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__8517\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__8514\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__8511\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__8506\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__8503\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__1580\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__1578\ : Span4Mux_h
    port map (
            O => \N__8486\,
            I => \N__8483\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__8483\,
            I => \uu2.mem0.N_10_0\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__8480\,
            I => \uu2.w_addr_displaying_4_rep1_3_cascade_\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__1574\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8468\
        );

    \I__1573\ : InMux
    port map (
            O => \N__8473\,
            I => \N__8468\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__8468\,
            I => \N__8463\
        );

    \I__1571\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8456\
        );

    \I__1570\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8456\
        );

    \I__1569\ : Span4Mux_h
    port map (
            O => \N__8463\,
            I => \N__8453\
        );

    \I__1568\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8448\
        );

    \I__1567\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8448\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__8456\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__8453\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__8448\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__1562\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8432\
        );

    \I__1561\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8432\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__8432\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__1559\ : InMux
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__8426\,
            I => \uu2.mem0.un1_segment4_0_i_i_1\
        );

    \I__1557\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__8420\,
            I => \uu2.mem0.un1_segment4_0_i_i_a5_0_0\
        );

    \I__1555\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8413\
        );

    \I__1554\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8410\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__8413\,
            I => \N__8403\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__8410\,
            I => \N__8400\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__8409\,
            I => \N__8393\
        );

    \I__1550\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8390\
        );

    \I__1549\ : InMux
    port map (
            O => \N__8407\,
            I => \N__8387\
        );

    \I__1548\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8384\
        );

    \I__1547\ : Span4Mux_h
    port map (
            O => \N__8403\,
            I => \N__8381\
        );

    \I__1546\ : Span4Mux_h
    port map (
            O => \N__8400\,
            I => \N__8378\
        );

    \I__1545\ : InMux
    port map (
            O => \N__8399\,
            I => \N__8375\
        );

    \I__1544\ : InMux
    port map (
            O => \N__8398\,
            I => \N__8366\
        );

    \I__1543\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8366\
        );

    \I__1542\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8366\
        );

    \I__1541\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8366\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__8390\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__8387\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__8384\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__8381\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__8378\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__8375\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__8366\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__8351\,
            I => \uu2.g1_0_1_cascade_\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__8348\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_50_cascade_\
        );

    \I__1531\ : InMux
    port map (
            O => \N__8345\,
            I => \N__8342\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__8342\,
            I => \uu2.g1_0_1\
        );

    \I__1529\ : InMux
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__8336\,
            I => \uu2.mem0.g0_0\
        );

    \I__1527\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8329\
        );

    \I__1526\ : InMux
    port map (
            O => \N__8332\,
            I => \N__8325\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__8329\,
            I => \N__8321\
        );

    \I__1524\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8318\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__8325\,
            I => \N__8315\
        );

    \I__1522\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8305\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__8321\,
            I => \N__8302\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__8318\,
            I => \N__8297\
        );

    \I__1519\ : Span4Mux_h
    port map (
            O => \N__8315\,
            I => \N__8297\
        );

    \I__1518\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8292\
        );

    \I__1517\ : InMux
    port map (
            O => \N__8313\,
            I => \N__8292\
        );

    \I__1516\ : InMux
    port map (
            O => \N__8312\,
            I => \N__8287\
        );

    \I__1515\ : InMux
    port map (
            O => \N__8311\,
            I => \N__8287\
        );

    \I__1514\ : InMux
    port map (
            O => \N__8310\,
            I => \N__8280\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8309\,
            I => \N__8280\
        );

    \I__1512\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8280\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__8305\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__8302\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1509\ : Odrv4
    port map (
            O => \N__8297\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__8292\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__8287\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__8280\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__8267\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__8264\,
            I => \N__8261\
        );

    \I__1503\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8258\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__8258\,
            I => \N__8255\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__8255\,
            I => \uu2.mem0.g1\
        );

    \I__1500\ : InMux
    port map (
            O => \N__8252\,
            I => \N__8243\
        );

    \I__1499\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8243\
        );

    \I__1498\ : InMux
    port map (
            O => \N__8250\,
            I => \N__8243\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__8243\,
            I => \uu2.N_10\
        );

    \I__1496\ : InMux
    port map (
            O => \N__8240\,
            I => \N__8237\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__8237\,
            I => \uu2.mem0.g1_1_1\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__8234\,
            I => \uu2.mem0.w_data_ns_1_1_0_3_cascade_\
        );

    \I__1493\ : InMux
    port map (
            O => \N__8231\,
            I => \N__8224\
        );

    \I__1492\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8224\
        );

    \I__1491\ : InMux
    port map (
            O => \N__8229\,
            I => \N__8221\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__8224\,
            I => \uu2.Z_decfrac106\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__8221\,
            I => \uu2.Z_decfrac106\
        );

    \I__1488\ : InMux
    port map (
            O => \N__8216\,
            I => \N__8213\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__8213\,
            I => \uu2.mem0.w_data_ns_1_0_0_1_3\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__8210\,
            I => \uu2.g0_1_0_0_1_cascade_\
        );

    \I__1485\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8201\
        );

    \I__1484\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8201\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__8201\,
            I => \uu2.g0_1_0_0\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1481\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__8192\,
            I => \uu2.g0_1_a5_0_0\
        );

    \I__1479\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__8186\,
            I => \N__8183\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__8183\,
            I => \uu2.g0_1_a5_1_0\
        );

    \I__1476\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8174\
        );

    \I__1475\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8174\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__8174\,
            I => \uu2.g1_1\
        );

    \I__1473\ : InMux
    port map (
            O => \N__8171\,
            I => \N__8168\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__8168\,
            I => \N__8162\
        );

    \I__1471\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8159\
        );

    \I__1470\ : InMux
    port map (
            O => \N__8166\,
            I => \N__8154\
        );

    \I__1469\ : InMux
    port map (
            O => \N__8165\,
            I => \N__8154\
        );

    \I__1468\ : Span4Mux_h
    port map (
            O => \N__8162\,
            I => \N__8151\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__8159\,
            I => \N__8148\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__8154\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__8151\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__8148\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1463\ : InMux
    port map (
            O => \N__8141\,
            I => \N__8128\
        );

    \I__1462\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8128\
        );

    \I__1461\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8128\
        );

    \I__1460\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8128\
        );

    \I__1459\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8125\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__8128\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__8125\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8116\
        );

    \I__1455\ : CascadeMux
    port map (
            O => \N__8119\,
            I => \N__8112\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__8116\,
            I => \N__8107\
        );

    \I__1453\ : InMux
    port map (
            O => \N__8115\,
            I => \N__8104\
        );

    \I__1452\ : InMux
    port map (
            O => \N__8112\,
            I => \N__8097\
        );

    \I__1451\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8097\
        );

    \I__1450\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8097\
        );

    \I__1449\ : Span4Mux_h
    port map (
            O => \N__8107\,
            I => \N__8092\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__8104\,
            I => \N__8092\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__8097\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__8092\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1445\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8082\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__8086\,
            I => \N__8078\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__8085\,
            I => \N__8075\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__8082\,
            I => \N__8071\
        );

    \I__1441\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8068\
        );

    \I__1440\ : InMux
    port map (
            O => \N__8078\,
            I => \N__8061\
        );

    \I__1439\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8061\
        );

    \I__1438\ : InMux
    port map (
            O => \N__8074\,
            I => \N__8061\
        );

    \I__1437\ : Span4Mux_v
    port map (
            O => \N__8071\,
            I => \N__8058\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__8068\,
            I => \N__8055\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__8061\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__8058\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__1433\ : Odrv4
    port map (
            O => \N__8055\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__8048\,
            I => \uu2.un2_w_addr_user_4_cascade_\
        );

    \I__1431\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8042\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__8042\,
            I => \N__8039\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__8039\,
            I => \uu2.un2_w_addr_user_5\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__8036\,
            I => \uu2.un448_ci_5_cascade_\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__8033\,
            I => \N__8028\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__8032\,
            I => \N__8025\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__8031\,
            I => \N__8022\
        );

    \I__1424\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8018\
        );

    \I__1423\ : InMux
    port map (
            O => \N__8025\,
            I => \N__8015\
        );

    \I__1422\ : InMux
    port map (
            O => \N__8022\,
            I => \N__8010\
        );

    \I__1421\ : InMux
    port map (
            O => \N__8021\,
            I => \N__8010\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__8018\,
            I => \N__8007\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__8015\,
            I => \N__8004\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__8010\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1417\ : Odrv4
    port map (
            O => \N__8007\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1416\ : Odrv12
    port map (
            O => \N__8004\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7997\,
            I => \N__7991\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7996\,
            I => \N__7991\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7991\,
            I => \N__7988\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__7988\,
            I => \N__7982\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7975\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7975\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7975\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__7982\,
            I => \uu2.un415_ci\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7975\,
            I => \uu2.un415_ci\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7963\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7954\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7968\,
            I => \N__7954\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7967\,
            I => \N__7954\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7954\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7963\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7954\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__7949\,
            I => \N__7946\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7943\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__7943\,
            I => \N__7940\
        );

    \I__1396\ : Odrv12
    port map (
            O => \N__7940\,
            I => \uu2.mem0.w_addr_4\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__7937\,
            I => \uu2.mem0.g0_8_0_cascade_\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7931\,
            I => \N__7924\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7930\,
            I => \N__7914\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7914\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7928\,
            I => \N__7914\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7927\,
            I => \N__7914\
        );

    \I__1388\ : Span4Mux_h
    port map (
            O => \N__7924\,
            I => \N__7911\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7923\,
            I => \N__7908\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7914\,
            I => \uu2.w_addr_userZ1Z_1\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__7911\,
            I => \uu2.w_addr_userZ1Z_1\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__7908\,
            I => \uu2.w_addr_userZ1Z_1\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__7901\,
            I => \uu2.o_adder_vbuf_w_addr_user_7_cascade_\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__7898\,
            I => \N__7895\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7892\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7892\,
            I => \N__7889\
        );

    \I__1379\ : Span4Mux_v
    port map (
            O => \N__7889\,
            I => \N__7886\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__7886\,
            I => \uu2.mem0.w_addr_7\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__7883\,
            I => \uu2.vbuf_w_addr_user.un459_ci_0_cascade_\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__7880\,
            I => \uu2.o_adder_vbuf_w_addr_user_8_cascade_\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7870\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7870\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7867\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7870\,
            I => \N__7864\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7867\,
            I => \uu2.un437_ci_3\
        );

    \I__1370\ : Odrv4
    port map (
            O => \N__7864\,
            I => \uu2.un437_ci_3\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7859\,
            I => \N__7855\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7858\,
            I => \N__7852\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7855\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7852\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7844\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7844\,
            I => vbuf_tx_data_0
        );

    \I__1363\ : InMux
    port map (
            O => \N__7841\,
            I => \N__7838\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7838\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7835\,
            I => \N__7832\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7832\,
            I => vbuf_tx_data_1
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7826\,
            I => \N__7823\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7823\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__7820\,
            I => \N__7817\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7814\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7814\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__7811\,
            I => \uu2.o_adder_vbuf_w_addr_user_3_cascade_\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7805\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7805\,
            I => \N__7800\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__7804\,
            I => \N__7796\
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__7803\,
            I => \N__7793\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__7800\,
            I => \N__7789\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7780\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7780\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7793\,
            I => \N__7780\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7792\,
            I => \N__7780\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__7789\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7780\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__7775\,
            I => \led_c_0_4_cascade_\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7772\,
            I => \N__7769\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7769\,
            I => \uu2.mem0.g1_0_0_0\
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__7766\,
            I => \N__7763\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7763\,
            I => \N__7760\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7760\,
            I => \uu2.mem0.g0_i_5_1_0\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7754\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7754\,
            I => \uu2.mem0.g2_0\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__7751\,
            I => \uu2.w_addr_displaying_4_rep1_8_cascade_\
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__7748\,
            I => \uu2.N_42_0_0_cascade_\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__7745\,
            I => \N__7742\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7742\,
            I => \N__7736\
        );

    \I__1329\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7736\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7736\,
            I => \N__7733\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__7733\,
            I => \uu2.N_1482_0_0\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__7730\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_34_cascade_\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__7727\,
            I => \uu2.mem0.un1_segment3_m6_0_0_0_0_cascade_\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7724\,
            I => \N__7721\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__7721\,
            I => \N__7718\
        );

    \I__1322\ : Span4Mux_h
    port map (
            O => \N__7718\,
            I => \N__7715\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__7715\,
            I => \uu2.mem0.w_data_3\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7712\,
            I => \N__7709\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7709\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_35\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7706\,
            I => \N__7703\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__7703\,
            I => \N__7700\
        );

    \I__1316\ : Odrv12
    port map (
            O => \N__7700\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_21\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7694\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7694\,
            I => \N__7691\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__7691\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_22\
        );

    \I__1312\ : InMux
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7685\,
            I => \N__7682\
        );

    \I__1310\ : Sp12to4
    port map (
            O => \N__7682\,
            I => \N__7679\
        );

    \I__1309\ : Odrv12
    port map (
            O => \N__7679\,
            I => \uu2.mem0.g0_i_a2_4\
        );

    \I__1308\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7673\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__7673\,
            I => \uu2.mem0.N_8_tz_0_0_1\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__7670\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_17_cascade_\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7667\,
            I => \N__7664\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__7664\,
            I => \N__7661\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__7661\,
            I => \uu2.mem0.w_data_5\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7658\,
            I => \N__7652\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7657\,
            I => \N__7652\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7652\,
            I => \uu2.Z_decfrac105_7_3\
        );

    \I__1299\ : CascadeMux
    port map (
            O => \N__7649\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_\
        );

    \I__1298\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__7643\,
            I => \N__7640\
        );

    \I__1296\ : Span4Mux_h
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__7637\,
            I => \uu2.mem0.w_data_0\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7634\,
            I => \N__7631\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__1292\ : Span4Mux_v
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__7625\,
            I => \uu2.mem0.w_data_2\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__7622\,
            I => \N__7619\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7619\,
            I => \N__7616\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__7616\,
            I => \uu2.un1_w_user_cr_0_0\
        );

    \I__1287\ : IoInMux
    port map (
            O => \N__7613\,
            I => \N__7610\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__7610\,
            I => \N__7606\
        );

    \I__1285\ : InMux
    port map (
            O => \N__7609\,
            I => \N__7603\
        );

    \I__1284\ : Span12Mux_s5_v
    port map (
            O => \N__7606\,
            I => \N__7598\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__7603\,
            I => \N__7598\
        );

    \I__1282\ : Odrv12
    port map (
            O => \N__7598\,
            I => \latticehx1k_pll_inst_PLLOUTCORE_i\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__7595\,
            I => \uu2.un1_w_user_cr_0_0_cascade_\
        );

    \I__1280\ : SRMux
    port map (
            O => \N__7592\,
            I => \N__7589\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__7589\,
            I => \N__7585\
        );

    \I__1278\ : CEMux
    port map (
            O => \N__7588\,
            I => \N__7582\
        );

    \I__1277\ : Span4Mux_v
    port map (
            O => \N__7585\,
            I => \N__7579\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__7582\,
            I => \N__7576\
        );

    \I__1275\ : Span4Mux_h
    port map (
            O => \N__7579\,
            I => \N__7571\
        );

    \I__1274\ : Span4Mux_v
    port map (
            O => \N__7576\,
            I => \N__7571\
        );

    \I__1273\ : Span4Mux_s2_h
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__7568\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1271\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7562\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__7562\,
            I => \resetGen.un3_reset_count_i_a3Z0Z_7\
        );

    \I__1269\ : InMux
    port map (
            O => \N__7559\,
            I => \N__7552\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7558\,
            I => \N__7552\
        );

    \I__1267\ : InMux
    port map (
            O => \N__7557\,
            I => \N__7549\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__7552\,
            I => \N__7546\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__7549\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1264\ : Odrv4
    port map (
            O => \N__7546\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__7541\,
            I => \N_87_cascade_\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7538\,
            I => \N__7534\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7537\,
            I => \N__7531\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__7534\,
            I => \N__7528\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__7531\,
            I => \N__7523\
        );

    \I__1258\ : Span4Mux_v
    port map (
            O => \N__7528\,
            I => \N__7523\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__7523\,
            I => \buart.Z_rx.N_91\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__7520\,
            I => \buart.Z_rx.N_91_cascade_\
        );

    \I__1255\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7514\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__7514\,
            I => \N__7508\
        );

    \I__1253\ : InMux
    port map (
            O => \N__7513\,
            I => \N__7505\
        );

    \I__1252\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7500\
        );

    \I__1251\ : InMux
    port map (
            O => \N__7511\,
            I => \N__7500\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__7508\,
            I => \buart.Z_rx.N_29_0_i_2\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__7505\,
            I => \buart.Z_rx.N_29_0_i_2\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__7500\,
            I => \buart.Z_rx.N_29_0_i_2\
        );

    \I__1247\ : InMux
    port map (
            O => \N__7493\,
            I => \N__7490\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__1245\ : Span4Mux_h
    port map (
            O => \N__7487\,
            I => \N__7484\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__7484\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__7481\,
            I => \buart.Z_rx.N_29_0_i_2_cascade_\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__7478\,
            I => \N__7475\
        );

    \I__1241\ : InMux
    port map (
            O => \N__7475\,
            I => \N__7471\
        );

    \I__1240\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7465\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__7471\,
            I => \N__7462\
        );

    \I__1238\ : InMux
    port map (
            O => \N__7470\,
            I => \N__7455\
        );

    \I__1237\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7455\
        );

    \I__1236\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7455\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__7465\,
            I => \N__7446\
        );

    \I__1234\ : Span4Mux_h
    port map (
            O => \N__7462\,
            I => \N__7446\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__7455\,
            I => \N__7446\
        );

    \I__1232\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7437\
        );

    \I__1231\ : InMux
    port map (
            O => \N__7453\,
            I => \N__7437\
        );

    \I__1230\ : Span4Mux_v
    port map (
            O => \N__7446\,
            I => \N__7434\
        );

    \I__1229\ : InMux
    port map (
            O => \N__7445\,
            I => \N__7425\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7425\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7443\,
            I => \N__7425\
        );

    \I__1226\ : InMux
    port map (
            O => \N__7442\,
            I => \N__7425\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__7437\,
            I => \buart.Z_rx.startbit\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__7434\,
            I => \buart.Z_rx.startbit\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__7425\,
            I => \buart.Z_rx.startbit\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__7418\,
            I => \N__7414\
        );

    \I__1221\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7411\
        );

    \I__1220\ : InMux
    port map (
            O => \N__7414\,
            I => \N__7406\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__7411\,
            I => \N__7403\
        );

    \I__1218\ : InMux
    port map (
            O => \N__7410\,
            I => \N__7398\
        );

    \I__1217\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7398\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__7406\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1215\ : Odrv4
    port map (
            O => \N__7403\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__7398\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1213\ : CEMux
    port map (
            O => \N__7391\,
            I => \N__7387\
        );

    \I__1212\ : CEMux
    port map (
            O => \N__7390\,
            I => \N__7384\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__7387\,
            I => \N__7380\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__7384\,
            I => \N__7377\
        );

    \I__1209\ : CEMux
    port map (
            O => \N__7383\,
            I => \N__7374\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__7380\,
            I => \N__7367\
        );

    \I__1207\ : Span4Mux_v
    port map (
            O => \N__7377\,
            I => \N__7367\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__7374\,
            I => \N__7367\
        );

    \I__1205\ : Span4Mux_v
    port map (
            O => \N__7367\,
            I => \N__7364\
        );

    \I__1204\ : Sp12to4
    port map (
            O => \N__7364\,
            I => \N__7361\
        );

    \I__1203\ : Odrv12
    port map (
            O => \N__7361\,
            I => \buart.Z_rx.bitcounte_0_i_2\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__7358\,
            I => \uu2.Z_decfrac105_7_3_cascade_\
        );

    \I__1201\ : InMux
    port map (
            O => \N__7355\,
            I => \N__7352\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__7352\,
            I => \N__7349\
        );

    \I__1199\ : Odrv12
    port map (
            O => \N__7349\,
            I => \uu2.mem0.w_data_6\
        );

    \I__1198\ : InMux
    port map (
            O => \N__7346\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__1197\ : InMux
    port map (
            O => \N__7343\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__1196\ : InMux
    port map (
            O => \N__7340\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__7337\,
            I => \N__7334\
        );

    \I__1194\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7331\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__7331\,
            I => \N__7328\
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__7328\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__7325\,
            I => \N__7322\
        );

    \I__1190\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7319\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__7319\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__1188\ : InMux
    port map (
            O => \N__7316\,
            I => \N__7313\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__7313\,
            I => \N__7310\
        );

    \I__1186\ : Span4Mux_h
    port map (
            O => \N__7310\,
            I => \N__7307\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__7307\,
            I => \uu2.mem0.w_data_7\
        );

    \I__1184\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7301\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__7301\,
            I => \N__7297\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__7300\,
            I => \N__7292\
        );

    \I__1181\ : Span4Mux_v
    port map (
            O => \N__7297\,
            I => \N__7289\
        );

    \I__1180\ : InMux
    port map (
            O => \N__7296\,
            I => \N__7282\
        );

    \I__1179\ : InMux
    port map (
            O => \N__7295\,
            I => \N__7282\
        );

    \I__1178\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7282\
        );

    \I__1177\ : Odrv4
    port map (
            O => \N__7289\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__7282\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__7277\,
            I => \buart.Z_rx.N_103_cascade_\
        );

    \I__1174\ : InMux
    port map (
            O => \N__7274\,
            I => \N__7271\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__7271\,
            I => \N__7268\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__7268\,
            I => \N__7265\
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__7265\,
            I => \uu2.r_data_wire_7\
        );

    \I__1170\ : InMux
    port map (
            O => \N__7262\,
            I => \N__7259\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__7259\,
            I => \N__7256\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__7256\,
            I => vbuf_tx_data_7
        );

    \I__1167\ : CEMux
    port map (
            O => \N__7253\,
            I => \N__7250\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__7250\,
            I => \N__7247\
        );

    \I__1165\ : Span4Mux_v
    port map (
            O => \N__7247\,
            I => \N__7243\
        );

    \I__1164\ : CEMux
    port map (
            O => \N__7246\,
            I => \N__7240\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__7243\,
            I => \uu2.vbuf_tx_data_rdy_0\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__7240\,
            I => \uu2.vbuf_tx_data_rdy_0\
        );

    \I__1161\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7232\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__7232\,
            I => vbuf_tx_data_3
        );

    \I__1159\ : InMux
    port map (
            O => \N__7229\,
            I => \N__7226\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__7226\,
            I => vbuf_tx_data_4
        );

    \I__1157\ : InMux
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__7220\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__7217\,
            I => \N__7214\
        );

    \I__1154\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7211\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__7211\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__1152\ : InMux
    port map (
            O => \N__7208\,
            I => \N__7205\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__7205\,
            I => vbuf_tx_data_2
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__7202\,
            I => \N__7199\
        );

    \I__1149\ : InMux
    port map (
            O => \N__7199\,
            I => \N__7196\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__7196\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__1147\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7190\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__7190\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__1145\ : IoInMux
    port map (
            O => \N__7187\,
            I => \N__7184\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__7184\,
            I => \N__7181\
        );

    \I__1143\ : IoSpan4Mux
    port map (
            O => \N__7181\,
            I => \N__7178\
        );

    \I__1142\ : Span4Mux_s3_h
    port map (
            O => \N__7178\,
            I => \N__7175\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__7175\,
            I => o_serial_data_c
        );

    \I__1140\ : InMux
    port map (
            O => \N__7172\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__7169\,
            I => \buart.Z_rx.ser_clk_cascade_\
        );

    \I__1138\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7163\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__7163\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__7160\,
            I => \N__7157\
        );

    \I__1135\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7152\
        );

    \I__1134\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7147\
        );

    \I__1133\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7147\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__7152\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__7147\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1130\ : InMux
    port map (
            O => \N__7142\,
            I => \N__7139\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__7139\,
            I => \N__7136\
        );

    \I__1128\ : Span4Mux_h
    port map (
            O => \N__7136\,
            I => \N__7133\
        );

    \I__1127\ : Span4Mux_v
    port map (
            O => \N__7133\,
            I => \N__7130\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__7130\,
            I => \uu2.r_data_wire_0\
        );

    \I__1125\ : InMux
    port map (
            O => \N__7127\,
            I => \N__7124\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__7124\,
            I => \N__7121\
        );

    \I__1123\ : Span4Mux_h
    port map (
            O => \N__7121\,
            I => \N__7118\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__7118\,
            I => \N__7115\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__7115\,
            I => \uu2.r_data_wire_1\
        );

    \I__1120\ : InMux
    port map (
            O => \N__7112\,
            I => \N__7109\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__7109\,
            I => \N__7106\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__7106\,
            I => \N__7103\
        );

    \I__1117\ : Span4Mux_v
    port map (
            O => \N__7103\,
            I => \N__7100\
        );

    \I__1116\ : Odrv4
    port map (
            O => \N__7100\,
            I => \uu2.r_data_wire_2\
        );

    \I__1115\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7094\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__7094\,
            I => \N__7091\
        );

    \I__1113\ : Span12Mux_s9_v
    port map (
            O => \N__7091\,
            I => \N__7088\
        );

    \I__1112\ : Odrv12
    port map (
            O => \N__7088\,
            I => \uu2.r_data_wire_3\
        );

    \I__1111\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7082\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__1109\ : Span4Mux_v
    port map (
            O => \N__7079\,
            I => \N__7076\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__7076\,
            I => \uu2.r_data_wire_4\
        );

    \I__1107\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7070\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__7070\,
            I => \N__7067\
        );

    \I__1105\ : Span4Mux_h
    port map (
            O => \N__7067\,
            I => \N__7064\
        );

    \I__1104\ : Span4Mux_v
    port map (
            O => \N__7064\,
            I => \N__7061\
        );

    \I__1103\ : Odrv4
    port map (
            O => \N__7061\,
            I => \uu2.r_data_wire_5\
        );

    \I__1102\ : InMux
    port map (
            O => \N__7058\,
            I => \N__7055\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__7055\,
            I => \N__7052\
        );

    \I__1100\ : Odrv4
    port map (
            O => \N__7052\,
            I => vbuf_tx_data_5
        );

    \I__1099\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7046\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__7046\,
            I => \N__7043\
        );

    \I__1097\ : Span12Mux_s9_h
    port map (
            O => \N__7043\,
            I => \N__7040\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__7040\,
            I => \uu2.r_data_wire_6\
        );

    \I__1095\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7034\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__7034\,
            I => vbuf_tx_data_6
        );

    \I__1093\ : InMux
    port map (
            O => \N__7031\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__1092\ : InMux
    port map (
            O => \N__7028\,
            I => \N__7025\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__7025\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__1089\ : InMux
    port map (
            O => \N__7019\,
            I => \N__7016\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__7016\,
            I => \N__7013\
        );

    \I__1087\ : Span4Mux_h
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__1086\ : Odrv4
    port map (
            O => \N__7010\,
            I => \uu2.mem0.g0_0_a3_0\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__7007\,
            I => \buart.Z_rx.startbit_cascade_\
        );

    \I__1084\ : InMux
    port map (
            O => \N__7004\,
            I => \N__6998\
        );

    \I__1083\ : InMux
    port map (
            O => \N__7003\,
            I => \N__6998\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__6998\,
            I => \N__6995\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__6995\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6992\,
            I => \N__6988\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6991\,
            I => \N__6985\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6988\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6985\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__6980\,
            I => \N__6977\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6970\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6970\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6967\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__6970\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6967\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__6962\,
            I => \N__6958\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__6961\,
            I => \N__6955\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6952\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6949\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6952\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__6949\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6939\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6934\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6934\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6939\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6934\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__6929\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__6926\,
            I => \N__6920\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6913\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6913\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6913\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6920\,
            I => \N__6910\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6913\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6910\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6905\,
            I => \N__6902\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6902\,
            I => \uu2.mem0.g0_i_5\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6899\,
            I => \N__6896\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6896\,
            I => \uu2.mem0.g0_i_6_1_0\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__6893\,
            I => \uu2.mem0.N_19_cascade_\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6890\,
            I => \N__6887\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6887\,
            I => \uu2.mem0.g0_i_6\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6881\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_53\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6878\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6875\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6872\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__6869\,
            I => \uu2.mem0.g2_1_0_0_cascade_\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6866\,
            I => \N__6863\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6863\,
            I => \uu2.mem0.g0_2_1\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__6860\,
            I => \uu2.mem0.g0_i_a2_3_cascade_\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6857\,
            I => \N__6854\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6854\,
            I => \uu2.mem0.w_data_displaying_2_0_0\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6848\,
            I => \uu2.mem0.g1_0_5\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6845\,
            I => \N__6842\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6842\,
            I => \uu2.mem0.N_10_0_0\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6839\,
            I => \N__6836\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6833\
        );

    \I__1027\ : Odrv4
    port map (
            O => \N__6833\,
            I => \uu2.mem0.g1_2\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__6830\,
            I => \N__6827\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6827\,
            I => \N__6824\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__6824\,
            I => \uu2.mem0.g1_1_sx\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6818\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6818\,
            I => \N__6815\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__6815\,
            I => \uu2.mem0.g1_0\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__6812\,
            I => \resetGen.N_104_cascade_\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6806\,
            I => \resetGen.N_84\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6803\,
            I => \N__6791\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6802\,
            I => \N__6791\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6801\,
            I => \N__6791\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6800\,
            I => \N__6791\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6791\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6779\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6787\,
            I => \N__6779\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6786\,
            I => \N__6779\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6779\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__6776\,
            I => \N__6773\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6769\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6766\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__6769\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6766\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6758\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6758\,
            I => \resetGen.N_86\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6755\,
            I => \N__6743\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6754\,
            I => \N__6743\
        );

    \I__999\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6743\
        );

    \I__998\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6743\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6743\,
            I => \resetGen.N_104\
        );

    \I__996\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6734\
        );

    \I__995\ : InMux
    port map (
            O => \N__6739\,
            I => \N__6734\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__6734\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__6731\,
            I => \resetGen.N_86_cascade_\
        );

    \I__992\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6724\
        );

    \I__991\ : CascadeMux
    port map (
            O => \N__6727\,
            I => \N__6720\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6724\,
            I => \N__6714\
        );

    \I__989\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6710\
        );

    \I__988\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6701\
        );

    \I__987\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6701\
        );

    \I__986\ : InMux
    port map (
            O => \N__6718\,
            I => \N__6701\
        );

    \I__985\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6701\
        );

    \I__984\ : Span4Mux_h
    port map (
            O => \N__6714\,
            I => \N__6698\
        );

    \I__983\ : InMux
    port map (
            O => \N__6713\,
            I => \N__6695\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__6710\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__6701\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__6698\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__6695\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__978\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__6683\,
            I => \Lab_UT.secuu0.un4_l_count_12\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__6680\,
            I => \N__6677\
        );

    \I__975\ : InMux
    port map (
            O => \N__6677\,
            I => \N__6674\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__6674\,
            I => \Lab_UT.secuu0.un87_ci\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__6671\,
            I => \Lab_UT.secuu0.un87_ci_cascade_\
        );

    \I__972\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6661\
        );

    \I__971\ : InMux
    port map (
            O => \N__6667\,
            I => \N__6661\
        );

    \I__970\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6658\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6661\,
            I => \Lab_UT.secuu0.l_countZ0Z_3\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__6658\,
            I => \Lab_UT.secuu0.l_countZ0Z_3\
        );

    \I__967\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6643\
        );

    \I__966\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6643\
        );

    \I__965\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6643\
        );

    \I__964\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6640\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6643\,
            I => \Lab_UT.secuu0.l_countZ0Z_2\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__6640\,
            I => \Lab_UT.secuu0.l_countZ0Z_2\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__6635\,
            I => \N__6629\
        );

    \I__960\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6625\
        );

    \I__959\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6618\
        );

    \I__958\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6618\
        );

    \I__957\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6618\
        );

    \I__956\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6615\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__6625\,
            I => \Lab_UT.secuu0.l_countZ0Z_0\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__6618\,
            I => \Lab_UT.secuu0.l_countZ0Z_0\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__6615\,
            I => \Lab_UT.secuu0.l_countZ0Z_0\
        );

    \I__952\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6602\
        );

    \I__951\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6595\
        );

    \I__950\ : InMux
    port map (
            O => \N__6606\,
            I => \N__6595\
        );

    \I__949\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6595\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__6602\,
            I => \N__6592\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__6595\,
            I => \Lab_UT.secuu0.l_countZ0Z_1\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__6592\,
            I => \Lab_UT.secuu0.l_countZ0Z_1\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__6587\,
            I => \Lab_UT.secuu0.un109_ci_cascade_\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__6584\,
            I => \N__6578\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__6583\,
            I => \N__6569\
        );

    \I__942\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6565\
        );

    \I__941\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6562\
        );

    \I__940\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6557\
        );

    \I__939\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6557\
        );

    \I__938\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6546\
        );

    \I__937\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6546\
        );

    \I__936\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6546\
        );

    \I__935\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6546\
        );

    \I__934\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6546\
        );

    \I__933\ : InMux
    port map (
            O => \N__6569\,
            I => \N__6541\
        );

    \I__932\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6541\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__6565\,
            I => \Lab_UT.secuu0.un153_ci\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__6562\,
            I => \Lab_UT.secuu0.un153_ci\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__6557\,
            I => \Lab_UT.secuu0.un153_ci\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__6546\,
            I => \Lab_UT.secuu0.un153_ci\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__6541\,
            I => \Lab_UT.secuu0.un153_ci\
        );

    \I__926\ : InMux
    port map (
            O => \N__6530\,
            I => \N__6524\
        );

    \I__925\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6524\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__6524\,
            I => \N__6521\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__6521\,
            I => \Lab_UT.secuu0.un131_ci_3\
        );

    \I__922\ : InMux
    port map (
            O => \N__6518\,
            I => \N__6514\
        );

    \I__921\ : InMux
    port map (
            O => \N__6517\,
            I => \N__6509\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__6514\,
            I => \N__6506\
        );

    \I__919\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6501\
        );

    \I__918\ : InMux
    port map (
            O => \N__6512\,
            I => \N__6501\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6509\,
            I => \N__6498\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__6506\,
            I => \Lab_UT.secuu0.l_countZ0Z_6\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__6501\,
            I => \Lab_UT.secuu0.l_countZ0Z_6\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__6498\,
            I => \Lab_UT.secuu0.l_countZ0Z_6\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__6491\,
            I => \N__6488\
        );

    \I__912\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6477\
        );

    \I__911\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6477\
        );

    \I__910\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6472\
        );

    \I__909\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6472\
        );

    \I__908\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6465\
        );

    \I__907\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6465\
        );

    \I__906\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6465\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__6477\,
            I => \N__6453\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__6472\,
            I => \N__6453\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__6465\,
            I => \N__6453\
        );

    \I__902\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6450\
        );

    \I__901\ : InMux
    port map (
            O => \N__6463\,
            I => \N__6441\
        );

    \I__900\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6441\
        );

    \I__899\ : InMux
    port map (
            O => \N__6461\,
            I => \N__6441\
        );

    \I__898\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6441\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__6453\,
            I => \Lab_UT.secuu0.un4_l_count_0\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__6450\,
            I => \Lab_UT.secuu0.un4_l_count_0\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__6441\,
            I => \Lab_UT.secuu0.un4_l_count_0\
        );

    \I__894\ : InMux
    port map (
            O => \N__6434\,
            I => \N__6431\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__6431\,
            I => \N__6428\
        );

    \I__892\ : Odrv12
    port map (
            O => \N__6428\,
            I => \Lab_UT.secuu0.un142_ci_0\
        );

    \I__891\ : InMux
    port map (
            O => \N__6425\,
            I => \N__6422\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__6422\,
            I => \N__6418\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__6421\,
            I => \N__6413\
        );

    \I__888\ : Span4Mux_h
    port map (
            O => \N__6418\,
            I => \N__6410\
        );

    \I__887\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6407\
        );

    \I__886\ : InMux
    port map (
            O => \N__6416\,
            I => \N__6402\
        );

    \I__885\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6402\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__6410\,
            I => \Lab_UT.secuu0.un109_ci\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__6407\,
            I => \Lab_UT.secuu0.un109_ci\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__6402\,
            I => \Lab_UT.secuu0.un109_ci\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__6395\,
            I => \N__6392\
        );

    \I__880\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6387\
        );

    \I__879\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6384\
        );

    \I__878\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6381\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__6387\,
            I => \Lab_UT.secuu0.l_countZ0Z_7\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__6384\,
            I => \Lab_UT.secuu0.l_countZ0Z_7\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__6381\,
            I => \Lab_UT.secuu0.l_countZ0Z_7\
        );

    \I__874\ : CEMux
    port map (
            O => \N__6374\,
            I => \N__6359\
        );

    \I__873\ : CEMux
    port map (
            O => \N__6373\,
            I => \N__6359\
        );

    \I__872\ : CEMux
    port map (
            O => \N__6372\,
            I => \N__6359\
        );

    \I__871\ : CEMux
    port map (
            O => \N__6371\,
            I => \N__6359\
        );

    \I__870\ : CEMux
    port map (
            O => \N__6370\,
            I => \N__6359\
        );

    \I__869\ : GlobalMux
    port map (
            O => \N__6359\,
            I => \N__6356\
        );

    \I__868\ : gio2CtrlBuf
    port map (
            O => \N__6356\,
            I => \Lab_UT.secuu0.un11_l_count_i_g\
        );

    \I__867\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6350\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__6350\,
            I => \Lab_UT.secuu0.un4_l_count_13\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__6347\,
            I => \Lab_UT.secuu0.un4_l_count_16_cascade_\
        );

    \I__864\ : InMux
    port map (
            O => \N__6344\,
            I => \N__6341\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__6338\,
            I => \Lab_UT.secuu0.un4_l_count_18\
        );

    \I__861\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6332\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__6332\,
            I => \Lab_UT.secuu0.delay_lineZ0Z_1\
        );

    \I__859\ : CascadeMux
    port map (
            O => \N__6329\,
            I => \Lab_UT.secuu0.un4_l_count_0_cascade_\
        );

    \I__858\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6322\
        );

    \I__857\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6319\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__6322\,
            I => \Lab_UT.secuu0.delay_lineZ0Z_0\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__6319\,
            I => \Lab_UT.secuu0.delay_lineZ0Z_0\
        );

    \I__854\ : IoInMux
    port map (
            O => \N__6314\,
            I => \N__6311\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__6311\,
            I => \N__6308\
        );

    \I__852\ : IoSpan4Mux
    port map (
            O => \N__6308\,
            I => \N__6305\
        );

    \I__851\ : Span4Mux_s0_h
    port map (
            O => \N__6305\,
            I => \N__6302\
        );

    \I__850\ : Span4Mux_h
    port map (
            O => \N__6302\,
            I => \N__6299\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__6299\,
            I => \Lab_UT.secuu0.un11_l_count_i\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__6296\,
            I => \N__6293\
        );

    \I__847\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6290\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__6290\,
            I => \Lab_UT.secuu0.un186_ci_0\
        );

    \I__845\ : InMux
    port map (
            O => \N__6287\,
            I => \N__6282\
        );

    \I__844\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6279\
        );

    \I__843\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6276\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__6282\,
            I => \Lab_UT.secuu0.l_countZ0Z_11\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__6279\,
            I => \Lab_UT.secuu0.l_countZ0Z_11\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__6276\,
            I => \Lab_UT.secuu0.l_countZ0Z_11\
        );

    \I__839\ : CascadeMux
    port map (
            O => \N__6269\,
            I => \N__6264\
        );

    \I__838\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6257\
        );

    \I__837\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6257\
        );

    \I__836\ : InMux
    port map (
            O => \N__6264\,
            I => \N__6257\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__6257\,
            I => \Lab_UT.secuu0.un241_ci_2\
        );

    \I__834\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6248\
        );

    \I__833\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6241\
        );

    \I__832\ : InMux
    port map (
            O => \N__6252\,
            I => \N__6241\
        );

    \I__831\ : InMux
    port map (
            O => \N__6251\,
            I => \N__6241\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__6248\,
            I => \N__6238\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__6241\,
            I => \Lab_UT.secuu0.l_countZ0Z_16\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__6238\,
            I => \Lab_UT.secuu0.l_countZ0Z_16\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__6233\,
            I => \Lab_UT.secuu0.un263_ci_cascade_\
        );

    \I__826\ : InMux
    port map (
            O => \N__6230\,
            I => \N__6226\
        );

    \I__825\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6223\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__6226\,
            I => \Lab_UT.secuu0.l_countZ0Z_18\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__6223\,
            I => \Lab_UT.secuu0.l_countZ0Z_18\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__6218\,
            I => \N__6214\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__6217\,
            I => \N__6209\
        );

    \I__820\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6205\
        );

    \I__819\ : InMux
    port map (
            O => \N__6213\,
            I => \N__6198\
        );

    \I__818\ : InMux
    port map (
            O => \N__6212\,
            I => \N__6198\
        );

    \I__817\ : InMux
    port map (
            O => \N__6209\,
            I => \N__6198\
        );

    \I__816\ : InMux
    port map (
            O => \N__6208\,
            I => \N__6195\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__6205\,
            I => \Lab_UT.secuu0.l_countZ0Z_9\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__6198\,
            I => \Lab_UT.secuu0.l_countZ0Z_9\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__6195\,
            I => \Lab_UT.secuu0.l_countZ0Z_9\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__6188\,
            I => \N__6183\
        );

    \I__811\ : InMux
    port map (
            O => \N__6187\,
            I => \N__6176\
        );

    \I__810\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6176\
        );

    \I__809\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6176\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__6176\,
            I => \Lab_UT.secuu0.l_countZ0Z_17\
        );

    \I__807\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6169\
        );

    \I__806\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6165\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__6169\,
            I => \N__6162\
        );

    \I__804\ : InMux
    port map (
            O => \N__6168\,
            I => \N__6159\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__6165\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__802\ : Odrv4
    port map (
            O => \N__6162\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__6159\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__6152\,
            I => \N__6148\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__6151\,
            I => \N__6145\
        );

    \I__798\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6140\
        );

    \I__797\ : InMux
    port map (
            O => \N__6145\,
            I => \N__6140\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__6140\,
            I => \uu2.vbuf_count.un372_ci_8_1\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__6137\,
            I => \N__6131\
        );

    \I__794\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6124\
        );

    \I__793\ : InMux
    port map (
            O => \N__6135\,
            I => \N__6124\
        );

    \I__792\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6124\
        );

    \I__791\ : InMux
    port map (
            O => \N__6131\,
            I => \N__6121\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__6124\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__6121\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__6116\,
            I => \uu2.vbuf_count.un372_ci_8_1_cascade_\
        );

    \I__787\ : InMux
    port map (
            O => \N__6113\,
            I => \N__6106\
        );

    \I__786\ : InMux
    port map (
            O => \N__6112\,
            I => \N__6106\
        );

    \I__785\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6103\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__6106\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__6103\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__782\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6094\
        );

    \I__781\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6089\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__6094\,
            I => \N__6086\
        );

    \I__779\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6081\
        );

    \I__778\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6081\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__6089\,
            I => \N__6078\
        );

    \I__776\ : Odrv4
    port map (
            O => \N__6086\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__6081\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__774\ : Odrv4
    port map (
            O => \N__6078\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__773\ : InMux
    port map (
            O => \N__6071\,
            I => \N__6068\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__6068\,
            I => \N__6061\
        );

    \I__771\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6054\
        );

    \I__770\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6054\
        );

    \I__769\ : InMux
    port map (
            O => \N__6065\,
            I => \N__6054\
        );

    \I__768\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6051\
        );

    \I__767\ : Odrv4
    port map (
            O => \N__6061\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__6054\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__6051\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__6044\,
            I => \N__6040\
        );

    \I__763\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6023\
        );

    \I__762\ : InMux
    port map (
            O => \N__6040\,
            I => \N__6023\
        );

    \I__761\ : InMux
    port map (
            O => \N__6039\,
            I => \N__6023\
        );

    \I__760\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6023\
        );

    \I__759\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6023\
        );

    \I__758\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6023\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__6023\,
            I => \N__6020\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__6020\,
            I => \uu2.un306_ci\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__6017\,
            I => \N__6010\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__6016\,
            I => \N__6006\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__6015\,
            I => \N__6003\
        );

    \I__752\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6000\
        );

    \I__751\ : InMux
    port map (
            O => \N__6013\,
            I => \N__5997\
        );

    \I__750\ : InMux
    port map (
            O => \N__6010\,
            I => \N__5988\
        );

    \I__749\ : InMux
    port map (
            O => \N__6009\,
            I => \N__5988\
        );

    \I__748\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5988\
        );

    \I__747\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5988\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__6000\,
            I => \N__5983\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5997\,
            I => \N__5983\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5988\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__743\ : Odrv12
    port map (
            O => \N__5983\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__5978\,
            I => \N__5972\
        );

    \I__741\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5965\
        );

    \I__740\ : InMux
    port map (
            O => \N__5976\,
            I => \N__5965\
        );

    \I__739\ : InMux
    port map (
            O => \N__5975\,
            I => \N__5965\
        );

    \I__738\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5962\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__5965\,
            I => \Lab_UT.secuu0.l_precountZ0Z_2\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5962\,
            I => \Lab_UT.secuu0.l_precountZ0Z_2\
        );

    \I__735\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5944\
        );

    \I__734\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5944\
        );

    \I__733\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5944\
        );

    \I__732\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5944\
        );

    \I__731\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5941\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__5944\,
            I => \Lab_UT.secuu0.l_precountZ0Z_1\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5941\,
            I => \Lab_UT.secuu0.l_precountZ0Z_1\
        );

    \I__728\ : InMux
    port map (
            O => \N__5936\,
            I => \N__5932\
        );

    \I__727\ : InMux
    port map (
            O => \N__5935\,
            I => \N__5928\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5932\,
            I => \N__5925\
        );

    \I__725\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5922\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5928\,
            I => \N__5917\
        );

    \I__723\ : Span4Mux_v
    port map (
            O => \N__5925\,
            I => \N__5917\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5922\,
            I => \Lab_UT.secuu0.l_countZ0Z_5\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__5917\,
            I => \Lab_UT.secuu0.l_countZ0Z_5\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__5912\,
            I => \N__5907\
        );

    \I__719\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5902\
        );

    \I__718\ : InMux
    port map (
            O => \N__5910\,
            I => \N__5902\
        );

    \I__717\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5899\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5902\,
            I => \Lab_UT.secuu0.l_precountZ0Z_3\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5899\,
            I => \Lab_UT.secuu0.l_precountZ0Z_3\
        );

    \I__714\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5887\
        );

    \I__713\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5887\
        );

    \I__712\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5884\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5887\,
            I => \Lab_UT.secuu0.l_countZ0Z_15\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5884\,
            I => \Lab_UT.secuu0.l_countZ0Z_15\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__5879\,
            I => \Lab_UT.secuu0.un4_l_count_11_cascade_\
        );

    \I__708\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5863\
        );

    \I__707\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5863\
        );

    \I__706\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5863\
        );

    \I__705\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5863\
        );

    \I__704\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5860\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5863\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5860\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__700\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5847\
        );

    \I__699\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5842\
        );

    \I__698\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5842\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5847\,
            I => \N__5839\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5842\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__695\ : Odrv12
    port map (
            O => \N__5839\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__5834\,
            I => \uu2.un3_r_clk_en_6_cascade_\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__5831\,
            I => \uu2_un3_r_clk_en_0_cascade_\
        );

    \I__692\ : CEMux
    port map (
            O => \N__5828\,
            I => \N__5824\
        );

    \I__691\ : SRMux
    port map (
            O => \N__5827\,
            I => \N__5821\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5824\,
            I => \N__5818\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5821\,
            I => \N__5809\
        );

    \I__688\ : Span4Mux_s3_h
    port map (
            O => \N__5818\,
            I => \N__5806\
        );

    \I__687\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5793\
        );

    \I__686\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5793\
        );

    \I__685\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5793\
        );

    \I__684\ : InMux
    port map (
            O => \N__5814\,
            I => \N__5793\
        );

    \I__683\ : InMux
    port map (
            O => \N__5813\,
            I => \N__5793\
        );

    \I__682\ : InMux
    port map (
            O => \N__5812\,
            I => \N__5793\
        );

    \I__681\ : Span4Mux_s3_h
    port map (
            O => \N__5809\,
            I => \N__5788\
        );

    \I__680\ : Span4Mux_h
    port map (
            O => \N__5806\,
            I => \N__5788\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5793\,
            I => \N__5785\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__5788\,
            I => \uu2.vbuf_tx_data_rdy\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__5785\,
            I => \uu2.vbuf_tx_data_rdy\
        );

    \I__676\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5777\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5777\,
            I => \uu2.un3_r_clk_en_0_0\
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__5774\,
            I => \N__5769\
        );

    \I__673\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5761\
        );

    \I__672\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5761\
        );

    \I__671\ : InMux
    port map (
            O => \N__5769\,
            I => \N__5761\
        );

    \I__670\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5758\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5761\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5758\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__5753\,
            I => \N__5749\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__5752\,
            I => \N__5746\
        );

    \I__665\ : InMux
    port map (
            O => \N__5749\,
            I => \N__5739\
        );

    \I__664\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5730\
        );

    \I__663\ : InMux
    port map (
            O => \N__5745\,
            I => \N__5730\
        );

    \I__662\ : InMux
    port map (
            O => \N__5744\,
            I => \N__5730\
        );

    \I__661\ : InMux
    port map (
            O => \N__5743\,
            I => \N__5730\
        );

    \I__660\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5727\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__5739\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5730\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5727\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__656\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5717\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__5717\,
            I => \uu2.un3_r_clk_en_7\
        );

    \I__654\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__5711\,
            I => \N__5708\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__5708\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__651\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5702\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5702\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__5699\,
            I => \uu2.un372_ci_cascade_\
        );

    \I__648\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5692\
        );

    \I__647\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5689\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__5692\,
            I => \uu2.l_countZ0Z_10\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__5689\,
            I => \uu2.l_countZ0Z_10\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__5684\,
            I => \uu2.un306_ci_cascade_\
        );

    \I__643\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__5678\,
            I => \uu2.un339_ci_0\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__640\ : InMux
    port map (
            O => \N__5672\,
            I => \N__5668\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__5671\,
            I => \N__5664\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__5668\,
            I => \N__5659\
        );

    \I__637\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5656\
        );

    \I__636\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5651\
        );

    \I__635\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5651\
        );

    \I__634\ : InMux
    port map (
            O => \N__5662\,
            I => \N__5648\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__5659\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__5656\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__5651\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__5648\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__628\ : InMux
    port map (
            O => \N__5636\,
            I => \N__5633\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5633\,
            I => \N__5627\
        );

    \I__626\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5624\
        );

    \I__625\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5621\
        );

    \I__624\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5618\
        );

    \I__623\ : Odrv4
    port map (
            O => \N__5627\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__5624\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__5621\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5618\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__5609\,
            I => \N__5604\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__5608\,
            I => \N__5601\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__5607\,
            I => \N__5598\
        );

    \I__616\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5595\
        );

    \I__615\ : InMux
    port map (
            O => \N__5601\,
            I => \N__5592\
        );

    \I__614\ : InMux
    port map (
            O => \N__5598\,
            I => \N__5589\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5595\,
            I => \N__5586\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__5592\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__5589\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__610\ : Odrv4
    port map (
            O => \N__5586\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__608\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__5573\,
            I => \N__5569\
        );

    \I__606\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5562\
        );

    \I__605\ : Span12Mux_s3_h
    port map (
            O => \N__5569\,
            I => \N__5559\
        );

    \I__604\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5556\
        );

    \I__603\ : InMux
    port map (
            O => \N__5567\,
            I => \N__5549\
        );

    \I__602\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5549\
        );

    \I__601\ : InMux
    port map (
            O => \N__5565\,
            I => \N__5549\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__5562\,
            I => \N__5546\
        );

    \I__599\ : Odrv12
    port map (
            O => \N__5559\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__5556\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__5549\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__596\ : Odrv4
    port map (
            O => \N__5546\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__595\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5526\
        );

    \I__594\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5526\
        );

    \I__593\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5526\
        );

    \I__592\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5521\
        );

    \I__591\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5521\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__5526\,
            I => \N__5518\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__5521\,
            I => \uu2.un415_ci_0\
        );

    \I__588\ : Odrv4
    port map (
            O => \N__5518\,
            I => \uu2.un415_ci_0\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__5513\,
            I => \uu2.vbuf_raddr.un459_ci_0_cascade_\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__5510\,
            I => \N__5507\
        );

    \I__585\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5503\
        );

    \I__584\ : InMux
    port map (
            O => \N__5506\,
            I => \N__5500\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__5503\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__5500\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__581\ : CascadeMux
    port map (
            O => \N__5495\,
            I => \N__5491\
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__5494\,
            I => \N__5488\
        );

    \I__579\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5483\
        );

    \I__578\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5476\
        );

    \I__577\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5476\
        );

    \I__576\ : InMux
    port map (
            O => \N__5486\,
            I => \N__5476\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__5483\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__5476\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__5471\,
            I => \N__5468\
        );

    \I__572\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5463\
        );

    \I__571\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5458\
        );

    \I__570\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5458\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__5463\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__5458\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__5453\,
            I => \N__5450\
        );

    \I__566\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5447\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__5447\,
            I => \N__5441\
        );

    \I__564\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5438\
        );

    \I__563\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5435\
        );

    \I__562\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5432\
        );

    \I__561\ : Odrv4
    port map (
            O => \N__5441\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__5438\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__5435\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__5432\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__556\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5416\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__5419\,
            I => \N__5412\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__5416\,
            I => \N__5407\
        );

    \I__553\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5404\
        );

    \I__552\ : InMux
    port map (
            O => \N__5412\,
            I => \N__5397\
        );

    \I__551\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5397\
        );

    \I__550\ : InMux
    port map (
            O => \N__5410\,
            I => \N__5397\
        );

    \I__549\ : Odrv4
    port map (
            O => \N__5407\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__5404\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__5397\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__5390\,
            I => \N__5387\
        );

    \I__545\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5381\
        );

    \I__544\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5381\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__5381\,
            I => \uu2.vbuf_raddr.un437_ci_3\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__5378\,
            I => \uu2.mem0.g0_0_a3_3_cascade_\
        );

    \I__541\ : InMux
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__5372\,
            I => \uu2.mem0.w_data_1\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__5369\,
            I => \uu2.mem0.g1_0_6_cascade_\
        );

    \I__538\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__5363\,
            I => \uu2.mem0.N_4_i\
        );

    \I__536\ : CascadeMux
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__535\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__5354\,
            I => \uu2.mem0.w_addr_6\
        );

    \I__533\ : InMux
    port map (
            O => \N__5351\,
            I => \N__5348\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__5348\,
            I => \uu2.mem0.N_14_0\
        );

    \I__531\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5342\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__5342\,
            I => \Lab_UT.secuu0.un208_ci_0\
        );

    \I__529\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5333\
        );

    \I__528\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5333\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__5333\,
            I => \Lab_UT.secuu0.l_countZ0Z_13\
        );

    \I__526\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5324\
        );

    \I__525\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5321\
        );

    \I__524\ : InMux
    port map (
            O => \N__5328\,
            I => \N__5318\
        );

    \I__523\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5315\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__5324\,
            I => \Lab_UT.secuu0.l_countZ0Z_10\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__5321\,
            I => \Lab_UT.secuu0.l_countZ0Z_10\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__5318\,
            I => \Lab_UT.secuu0.l_countZ0Z_10\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__5315\,
            I => \Lab_UT.secuu0.l_countZ0Z_10\
        );

    \I__518\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5294\
        );

    \I__517\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5294\
        );

    \I__516\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5294\
        );

    \I__515\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5287\
        );

    \I__514\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5287\
        );

    \I__513\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5287\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__5294\,
            I => \Lab_UT.secuu0.l_countZ0Z_8\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__5287\,
            I => \Lab_UT.secuu0.l_countZ0Z_8\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__5282\,
            I => \N__5279\
        );

    \I__509\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__5276\,
            I => \uu2.mem0.w_addr_8\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__506\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__5267\,
            I => \uu2.mem0.w_addr_1\
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__5264\,
            I => \N__5261\
        );

    \I__503\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__501\ : Odrv4
    port map (
            O => \N__5255\,
            I => \uu2.mem0.w_addr_2\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__499\ : InMux
    port map (
            O => \N__5249\,
            I => \N__5246\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__5246\,
            I => \uu2.mem0.w_addr_5\
        );

    \I__497\ : InMux
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__5240\,
            I => \uu2.mem0.w_data_4\
        );

    \I__495\ : CascadeMux
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__494\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5231\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__5231\,
            I => \uu2.mem0.w_addr_3\
        );

    \I__492\ : CascadeMux
    port map (
            O => \N__5228\,
            I => \Lab_UT.secuu0.un230_ci_1_cascade_\
        );

    \I__491\ : CascadeMux
    port map (
            O => \N__5225\,
            I => \N__5219\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__5224\,
            I => \N__5216\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__5223\,
            I => \N__5211\
        );

    \I__488\ : InMux
    port map (
            O => \N__5222\,
            I => \N__5208\
        );

    \I__487\ : InMux
    port map (
            O => \N__5219\,
            I => \N__5197\
        );

    \I__486\ : InMux
    port map (
            O => \N__5216\,
            I => \N__5197\
        );

    \I__485\ : InMux
    port map (
            O => \N__5215\,
            I => \N__5197\
        );

    \I__484\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5197\
        );

    \I__483\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5197\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__5208\,
            I => \N__5194\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__5197\,
            I => \Lab_UT.secuu0.l_precountZ0Z_0\
        );

    \I__480\ : Odrv4
    port map (
            O => \N__5194\,
            I => \Lab_UT.secuu0.l_precountZ0Z_0\
        );

    \I__479\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5185\
        );

    \I__478\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5182\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__5185\,
            I => \N__5178\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__5182\,
            I => \N__5174\
        );

    \I__475\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5171\
        );

    \I__474\ : Span4Mux_s3_h
    port map (
            O => \N__5178\,
            I => \N__5168\
        );

    \I__473\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5165\
        );

    \I__472\ : Odrv4
    port map (
            O => \N__5174\,
            I => \Lab_UT.secuu0.l_countZ0Z_4\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__5171\,
            I => \Lab_UT.secuu0.l_countZ0Z_4\
        );

    \I__470\ : Odrv4
    port map (
            O => \N__5168\,
            I => \Lab_UT.secuu0.l_countZ0Z_4\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__5165\,
            I => \Lab_UT.secuu0.l_countZ0Z_4\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__5156\,
            I => \Lab_UT.secuu0.un4_l_count_14_cascade_\
        );

    \I__467\ : InMux
    port map (
            O => \N__5153\,
            I => \N__5146\
        );

    \I__466\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5146\
        );

    \I__465\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5143\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__5146\,
            I => \Lab_UT.secuu0.un4_l_count_0_8\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__5143\,
            I => \Lab_UT.secuu0.un4_l_count_0_8\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__5138\,
            I => \Lab_UT.secuu0.un4_l_count_0_8_cascade_\
        );

    \I__461\ : CascadeMux
    port map (
            O => \N__5135\,
            I => \N__5129\
        );

    \I__460\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5124\
        );

    \I__459\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5124\
        );

    \I__458\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5119\
        );

    \I__457\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5119\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__5124\,
            I => \Lab_UT.secuu0.l_countZ0Z_14\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__5119\,
            I => \Lab_UT.secuu0.l_countZ0Z_14\
        );

    \I__454\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5106\
        );

    \I__453\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5106\
        );

    \I__452\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5101\
        );

    \I__451\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5101\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__5106\,
            I => \Lab_UT.secuu0.un197_ci_9\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__5101\,
            I => \Lab_UT.secuu0.un197_ci_9\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__447\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5088\
        );

    \I__446\ : InMux
    port map (
            O => \N__5092\,
            I => \N__5085\
        );

    \I__445\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5082\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__5088\,
            I => \Lab_UT.secuu0.l_countZ0Z_12\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__5085\,
            I => \Lab_UT.secuu0.l_countZ0Z_12\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__5082\,
            I => \Lab_UT.secuu0.l_countZ0Z_12\
        );

    \I__441\ : CascadeMux
    port map (
            O => \N__5075\,
            I => \Lab_UT.secuu0.un197_ci_9_cascade_\
        );

    \I__440\ : IoInMux
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__5069\,
            I => \resetGen.rst_isoZ0\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__5066\,
            I => \Lab_UT.secuu0.un131_ci_3_cascade_\
        );

    \I__437\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N__5057\
        );

    \I__435\ : Odrv4
    port map (
            O => \N__5057\,
            I => \uart_RXD\
        );

    \I__434\ : IoInMux
    port map (
            O => \N__5054\,
            I => \N__5051\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__5051\,
            I => \N__5048\
        );

    \I__432\ : IoSpan4Mux
    port map (
            O => \N__5048\,
            I => \N__5045\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__5045\,
            I => clk_in_c
        );

    \INVuu2.w_addr_displaying_fast_5C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_5C_net\,
            I => \N__13408\
        );

    \INVuu2.w_addr_displaying_8C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_8C_net\,
            I => \N__13396\
        );

    \INVuu2.w_addr_displaying_fast_1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_1C_net\,
            I => \N__13401\
        );

    \INVuu2.w_addr_displaying_fast_0C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_0C_net\,
            I => \N__13407\
        );

    \INVuu2.w_addr_displaying_fast_6C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_6C_net\,
            I => \N__13413\
        );

    \INVuu2.w_addr_user_0C\ : INV
    port map (
            O => \INVuu2.w_addr_user_0C_net\,
            I => \N__13430\
        );

    \INVuu2.w_addr_displaying_3_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_3_rep1C_net\,
            I => \N__13390\
        );

    \INVuu2.w_addr_displaying_0_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_0_rep1C_net\,
            I => \N__13395\
        );

    \INVuu2.w_addr_displaying_2_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_2_rep1C_net\,
            I => \N__13400\
        );

    \INVuu2.w_addr_displaying_5_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_5_rep1C_net\,
            I => \N__13406\
        );

    \INVuu2.w_addr_user_5C\ : INV
    port map (
            O => \INVuu2.w_addr_user_5C_net\,
            I => \N__13412\
        );

    \INVuu2.w_addr_user_7C\ : INV
    port map (
            O => \INVuu2.w_addr_user_7C_net\,
            I => \N__13417\
        );

    \INVuu2.w_addr_user_2C\ : INV
    port map (
            O => \INVuu2.w_addr_user_2C_net\,
            I => \N__13424\
        );

    \INVuu2.w_addr_displaying_8_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_8_rep1C_net\,
            I => \N__13383\
        );

    \INVuu2.w_addr_displaying_5C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_5C_net\,
            I => \N__13397\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_12_0_\
        );

    \resetGen.rst_iso_RNIEOGF\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5072\,
            GLOBALBUFFEROUTPUT => \resetGen_rst_iso_g\
        );

    \Lab_UT.secuu0.delay_line_RNILBAI7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6314\,
            GLOBALBUFFEROUTPUT => \Lab_UT.secuu0.un11_l_count_i_g\
        );

    \latticehx1k_pll_inst.PLLOUTCORE_derived_clock_RNIALC1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7613\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \resetGen.rst_iso_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6728\,
            lcout => \resetGen.rst_isoZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_5_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__6425\,
            in1 => \N__5188\,
            in2 => \_gnd_net_\,
            in3 => \N__5935\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13432\,
            ce => \N__6370\,
            sr => \N__12307\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_3_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5931\,
            in2 => \_gnd_net_\,
            in3 => \N__5189\,
            lcout => \Lab_UT.secuu0.un131_ci_3\,
            ltout => \Lab_UT.secuu0.un131_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_7__un142_ci_0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6518\,
            in2 => \N__5066\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.secuu0.un142_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_0_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5063\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13404\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.sec_clk_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6464\,
            in2 => \_gnd_net_\,
            in3 => \N__13107\,
            lcout => \Lab_UT_l_oneSecPluse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13429\,
            ce => 'H',
            sr => \N__12311\
        );

    \Lab_UT.secuu0.delay_line_1_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6326\,
            lcout => \Lab_UT.secuu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13429\,
            ce => 'H',
            sr => \N__12311\
        );

    \Lab_UT.secuu0.l_precount_0_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5214\,
            lcout => \Lab_UT.secuu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13429\,
            ce => 'H',
            sr => \N__12311\
        );

    \Lab_UT.secuu0.l_precount_3_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__5977\,
            in1 => \N__5911\,
            in2 => \N__5225\,
            in3 => \N__5957\,
            lcout => \Lab_UT.secuu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13429\,
            ce => 'H',
            sr => \N__12311\
        );

    \Lab_UT.secuu0.l_precount_2_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__5976\,
            in1 => \_gnd_net_\,
            in2 => \N__5224\,
            in3 => \N__5956\,
            lcout => \Lab_UT.secuu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13429\,
            ce => 'H',
            sr => \N__12311\
        );

    \Lab_UT.secuu0.l_precount_1_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__5955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5215\,
            lcout => \Lab_UT.secuu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13429\,
            ce => 'H',
            sr => \N__12311\
        );

    \Lab_UT.secuu0.delay_line_0_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5975\,
            in1 => \N__5910\,
            in2 => \N__5223\,
            in3 => \N__5954\,
            lcout => \Lab_UT.secuu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13429\,
            ce => 'H',
            sr => \N__12311\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_13__un208_ci_0_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5111\,
            in2 => \_gnd_net_\,
            in3 => \N__5092\,
            lcout => \Lab_UT.secuu0.un208_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_11__un186_ci_0_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5305\,
            in1 => \N__6212\,
            in2 => \_gnd_net_\,
            in3 => \N__5329\,
            lcout => \Lab_UT.secuu0.un186_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_12__un197_ci_9_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6286\,
            in1 => \N__5328\,
            in2 => \N__6217\,
            in3 => \N__5304\,
            lcout => \Lab_UT.secuu0.un197_ci_9\,
            ltout => \Lab_UT.secuu0.un197_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_16__un241_ci_2_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5893\,
            in1 => \N__5133\,
            in2 => \N__5075\,
            in3 => \N__5152\,
            lcout => \Lab_UT.secuu0.un241_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_9_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__6213\,
            in1 => \N__6582\,
            in2 => \_gnd_net_\,
            in3 => \N__5306\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13427\,
            ce => \N__6372\,
            sr => \N__12309\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_15__un230_ci_1_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5112\,
            in1 => \N__5134\,
            in2 => \_gnd_net_\,
            in3 => \N__5153\,
            lcout => OPEN,
            ltout => \Lab_UT.secuu0.un230_ci_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_15_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__6581\,
            in1 => \N__6485\,
            in2 => \N__5228\,
            in3 => \N__5894\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13427\,
            ce => \N__6372\,
            sr => \N__12309\
        );

    \Lab_UT.secuu0.l_count_4_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6486\,
            in1 => \N__6417\,
            in2 => \_gnd_net_\,
            in3 => \N__5181\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13427\,
            ce => \N__6372\,
            sr => \N__12309\
        );

    \Lab_UT.secuu0.l_count_RNI0S951_2_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5327\,
            in1 => \N__5301\,
            in2 => \N__5135\,
            in3 => \N__6650\,
            lcout => OPEN,
            ltout => \Lab_UT.secuu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_RNI20OC2_4_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5222\,
            in1 => \N__5177\,
            in2 => \N__5156\,
            in3 => \N__5151\,
            lcout => \Lab_UT.secuu0.un4_l_count_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_RNIFM2M_13_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5338\,
            in2 => \_gnd_net_\,
            in3 => \N__5091\,
            lcout => \Lab_UT.secuu0.un4_l_count_0_8\,
            ltout => \Lab_UT.secuu0.un4_l_count_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_14_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__5114\,
            in1 => \N__6575\,
            in2 => \N__5138\,
            in3 => \N__5132\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13422\,
            ce => \N__6371\,
            sr => \N__12308\
        );

    \Lab_UT.secuu0.l_count_12_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__6573\,
            in1 => \N__6487\,
            in2 => \N__5096\,
            in3 => \N__5113\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13422\,
            ce => \N__6371\,
            sr => \N__12308\
        );

    \Lab_UT.secuu0.l_count_13_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__5339\,
            in1 => \N__5345\,
            in2 => \N__6491\,
            in3 => \N__6574\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13422\,
            ce => \N__6371\,
            sr => \N__12308\
        );

    \Lab_UT.secuu0.l_count_10_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__6576\,
            in1 => \N__5330\,
            in2 => \N__6218\,
            in3 => \N__5302\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13422\,
            ce => \N__6371\,
            sr => \N__12308\
        );

    \Lab_UT.secuu0.l_count_8_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__5303\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6572\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13422\,
            ce => \N__6371\,
            sr => \N__12308\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11248\,
            in1 => \N__8171\,
            in2 => \_gnd_net_\,
            in3 => \N__9967\,
            lcout => \uu2.mem0.w_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7934\,
            in1 => \N__11249\,
            in2 => \_gnd_net_\,
            in3 => \N__11694\,
            lcout => \uu2.mem0.w_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11245\,
            in1 => \N__8120\,
            in2 => \_gnd_net_\,
            in3 => \N__11596\,
            lcout => \uu2.mem0.w_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__11247\,
            in1 => \_gnd_net_\,
            in2 => \N__8033\,
            in3 => \N__11872\,
            lcout => \uu2.mem0.w_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__10967\,
            in1 => \N__6857\,
            in2 => \_gnd_net_\,
            in3 => \N__11250\,
            lcout => \uu2.mem0.w_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11246\,
            in1 => \N__7808\,
            in2 => \_gnd_net_\,
            in3 => \N__12079\,
            lcout => \uu2.mem0.w_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_23_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6890\,
            in1 => \N__5351\,
            in2 => \N__7022\,
            in3 => \N__6905\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_0_a3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__6821\,
            in1 => \N__6866\,
            in2 => \N__5378\,
            in3 => \N__5366\,
            lcout => \uu2.mem0.w_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_31_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6884\,
            in2 => \_gnd_net_\,
            in3 => \N__6851\,
            lcout => OPEN,
            ltout => \uu2.mem0.g1_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_19_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010001000100"
        )
    port map (
            in0 => \N__6839\,
            in1 => \N__11251\,
            in2 => \N__5369\,
            in3 => \N__9707\,
            lcout => \uu2.mem0.N_4_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11252\,
            in1 => \N__8087\,
            in2 => \_gnd_net_\,
            in3 => \N__9865\,
            lcout => \uu2.mem0.w_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6713\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13410\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_36_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001000"
        )
    port map (
            in0 => \N__12077\,
            in1 => \N__8333\,
            in2 => \N__11597\,
            in3 => \N__8549\,
            lcout => \uu2.mem0.N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_3_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__5632\,
            in1 => \N__5667\,
            in2 => \N__5607\,
            in3 => \N__5568\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13405\,
            ce => \N__7246\,
            sr => \N__12298\
        );

    \uu2.r_addr_esr_6_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__5446\,
            in1 => \N__5415\,
            in2 => \N__5494\,
            in3 => \N__5535\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13405\,
            ce => \N__7246\,
            sr => \N__12298\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un459_ci_0_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5466\,
            in2 => \_gnd_net_\,
            in3 => \N__5486\,
            lcout => OPEN,
            ltout => \uu2.vbuf_raddr.un459_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_8_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__5506\,
            in1 => \N__5386\,
            in2 => \N__5513\,
            in3 => \N__5536\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13405\,
            ce => \N__7246\,
            sr => \N__12298\
        );

    \uu2.r_addr_esr_7_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__5537\,
            in1 => \N__5467\,
            in2 => \N__5390\,
            in3 => \N__5487\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13405\,
            ce => \N__7246\,
            sr => \N__12298\
        );

    \uu2.r_addr_2_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__5815\,
            in1 => \N__5631\,
            in2 => \N__5671\,
            in3 => \N__5567\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13398\,
            ce => 'H',
            sr => \N__12322\
        );

    \uu2.r_addr_1_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__5566\,
            in1 => \N__5663\,
            in2 => \_gnd_net_\,
            in3 => \N__5816\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13398\,
            ce => 'H',
            sr => \N__12322\
        );

    \uu2.r_addr_0_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__5813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5565\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13398\,
            ce => 'H',
            sr => \N__12322\
        );

    \uu2.l_count_RNI88MU5_4_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12321\,
            in2 => \_gnd_net_\,
            in3 => \N__5812\,
            lcout => \uu2.vbuf_tx_data_rdy_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_4_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__5814\,
            in1 => \N__5411\,
            in2 => \_gnd_net_\,
            in3 => \N__5533\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13398\,
            ce => 'H',
            sr => \N__12322\
        );

    \uu2.r_addr_5_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__5534\,
            in1 => \N__5445\,
            in2 => \N__5419\,
            in3 => \N__5817\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13398\,
            ce => 'H',
            sr => \N__12322\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un437_ci_3_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5444\,
            in2 => \_gnd_net_\,
            in3 => \N__5410\,
            lcout => \uu2.vbuf_raddr.un437_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_1_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5745\,
            in2 => \_gnd_net_\,
            in3 => \N__5874\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13393\,
            ce => 'H',
            sr => \N__12299\
        );

    \uu2.l_count_3_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__5876\,
            in1 => \N__5773\,
            in2 => \N__5752\,
            in3 => \N__5851\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13393\,
            ce => 'H',
            sr => \N__12299\
        );

    \uu2.l_count_2_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__5772\,
            in1 => \N__10476\,
            in2 => \N__5753\,
            in3 => \N__5875\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13393\,
            ce => 'H',
            sr => \N__12299\
        );

    \uu2.l_count_0_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__5744\,
            in1 => \_gnd_net_\,
            in2 => \N__10506\,
            in3 => \_gnd_net_\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13393\,
            ce => 'H',
            sr => \N__12299\
        );

    \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5850\,
            in1 => \N__5743\,
            in2 => \N__5774\,
            in3 => \N__5873\,
            lcout => \uu2.un306_ci\,
            ltout => \uu2.un306_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_7_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__10472\,
            in1 => \N__5681\,
            in2 => \N__5684\,
            in3 => \N__6172\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13393\,
            ce => 'H',
            sr => \N__12299\
        );

    \uu2.vbuf_count.counter_gen_label_7__un339_ci_0_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6014\,
            in1 => \N__6098\,
            in2 => \_gnd_net_\,
            in3 => \N__6071\,
            lcout => \uu2.un339_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un415_ci_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5662\,
            in1 => \N__5630\,
            in2 => \N__5609\,
            in3 => \N__5572\,
            lcout => \uu2.un415_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_6_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__10286\,
            in1 => \N__5714\,
            in2 => \N__10507\,
            in3 => \N__7058\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13388\,
            ce => \N__8588\,
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNICDGK1_3_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__6168\,
            in1 => \N__5872\,
            in2 => \N__5855\,
            in3 => \N__6111\,
            lcout => OPEN,
            ltout => \uu2.un3_r_clk_en_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI0NA44_4_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6013\,
            in1 => \N__5720\,
            in2 => \N__5834\,
            in3 => \N__5780\,
            lcout => uu2_un3_r_clk_en_0,
            ltout => \uu2_un3_r_clk_en_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIQF5F5_4_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5831\,
            in3 => \N__10285\,
            lcout => \uu2.vbuf_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI2U5E_10_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5695\,
            in2 => \_gnd_net_\,
            in3 => \N__6064\,
            lcout => \uu2.un3_r_clk_en_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI89GK1_2_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6097\,
            in1 => \N__5768\,
            in2 => \N__6137\,
            in3 => \N__5742\,
            lcout => \uu2.un3_r_clk_en_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_7_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__10287\,
            in1 => \N__5705\,
            in2 => \N__10508\,
            in3 => \N__7037\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13388\,
            ce => \N__8588\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_8_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__7262\,
            in1 => \N__10477\,
            in2 => \_gnd_net_\,
            in3 => \N__10288\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13388\,
            ce => \N__8588\,
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_10__un372_ci_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6036\,
            in1 => \N__6134\,
            in2 => \N__6151\,
            in3 => \N__6112\,
            lcout => OPEN,
            ltout => \uu2.un372_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_10_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__10469\,
            in1 => \_gnd_net_\,
            in2 => \N__5699\,
            in3 => \N__5696\,
            lcout => \uu2.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13384\,
            ce => 'H',
            sr => \N__12301\
        );

    \uu2.l_count_8_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__6037\,
            in1 => \_gnd_net_\,
            in2 => \N__6152\,
            in3 => \N__6135\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13384\,
            ce => 'H',
            sr => \N__12301\
        );

    \uu2.vbuf_count.counter_gen_label_10__un372_ci_8_1_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6092\,
            in1 => \N__6173\,
            in2 => \N__6015\,
            in3 => \N__6065\,
            lcout => \uu2.vbuf_count.un372_ci_8_1\,
            ltout => \uu2.vbuf_count.un372_ci_8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_9_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__6039\,
            in1 => \N__6136\,
            in2 => \N__6116\,
            in3 => \N__6113\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13384\,
            ce => 'H',
            sr => \N__12301\
        );

    \uu2.l_count_6_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__6093\,
            in1 => \N__6043\,
            in2 => \N__6017\,
            in3 => \N__6067\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13384\,
            ce => 'H',
            sr => \N__12301\
        );

    \uu2.l_count_5_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__6066\,
            in1 => \N__6009\,
            in2 => \N__6044\,
            in3 => \N__10471\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13384\,
            ce => 'H',
            sr => \N__12301\
        );

    \uu2.l_count_4_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000010100"
        )
    port map (
            in0 => \N__10470\,
            in1 => \N__6038\,
            in2 => \N__6016\,
            in3 => \_gnd_net_\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13384\,
            ce => 'H',
            sr => \N__12301\
        );

    \Lab_UT.secuu0.l_count_RNI24E71_11_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__6254\,
            in1 => \N__6628\,
            in2 => \N__5978\,
            in3 => \N__6285\,
            lcout => \Lab_UT.secuu0.un4_l_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_RNI8TM21_5_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5953\,
            in1 => \N__5936\,
            in2 => \N__5912\,
            in3 => \N__6608\,
            lcout => OPEN,
            ltout => \Lab_UT.secuu0.un4_l_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_RNI9GD02_18_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6229\,
            in1 => \N__5892\,
            in2 => \N__5879\,
            in3 => \N__6517\,
            lcout => OPEN,
            ltout => \Lab_UT.secuu0.un4_l_count_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_RNI82GM6_3_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6353\,
            in1 => \N__6686\,
            in2 => \N__6347\,
            in3 => \N__6344\,
            lcout => \Lab_UT.secuu0.un4_l_count_0\,
            ltout => \Lab_UT.secuu0.un4_l_count_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.delay_line_RNILBAI7_1_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6335\,
            in2 => \N__6329\,
            in3 => \N__6325\,
            lcout => \Lab_UT.secuu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_0_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6460\,
            in2 => \_gnd_net_\,
            in3 => \N__6634\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13423\,
            ce => \N__6374\,
            sr => \N__12312\
        );

    \Lab_UT.secuu0.l_count_11_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__6461\,
            in1 => \N__6577\,
            in2 => \N__6296\,
            in3 => \N__6287\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13423\,
            ce => \N__6374\,
            sr => \N__12312\
        );

    \Lab_UT.secuu0.l_count_16_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__6267\,
            in1 => \N__6462\,
            in2 => \N__6584\,
            in3 => \N__6252\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13423\,
            ce => \N__6374\,
            sr => \N__12312\
        );

    \Lab_UT.secuu0.l_count_17_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__6253\,
            in1 => \N__6268\,
            in2 => \N__6583\,
            in3 => \N__6187\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13423\,
            ce => \N__6374\,
            sr => \N__12312\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_18__un263_ci_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6186\,
            in1 => \N__6568\,
            in2 => \N__6269\,
            in3 => \N__6251\,
            lcout => OPEN,
            ltout => \Lab_UT.secuu0.un263_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_18_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__6463\,
            in1 => \_gnd_net_\,
            in2 => \N__6233\,
            in3 => \N__6230\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13423\,
            ce => \N__6374\,
            sr => \N__12312\
        );

    \Lab_UT.secuu0.l_count_RNIRDS11_3_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6208\,
            in1 => \N__6666\,
            in2 => \N__6188\,
            in3 => \N__6390\,
            lcout => \Lab_UT.secuu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_3_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__6668\,
            in1 => \N__6484\,
            in2 => \N__6680\,
            in3 => \N__6653\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13416\,
            ce => \N__6373\,
            sr => \N__12310\
        );

    \Lab_UT.secuu0.l_count_1_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__6607\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6633\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13416\,
            ce => \N__6373\,
            sr => \N__12310\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_1_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6632\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6606\,
            lcout => \Lab_UT.secuu0.un87_ci\,
            ltout => \Lab_UT.secuu0.un87_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_2_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__6652\,
            in1 => \_gnd_net_\,
            in2 => \N__6671\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13416\,
            ce => \N__6373\,
            sr => \N__12310\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_6_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6667\,
            in1 => \N__6651\,
            in2 => \N__6635\,
            in3 => \N__6605\,
            lcout => \Lab_UT.secuu0.un109_ci\,
            ltout => \Lab_UT.secuu0.un109_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_8_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6529\,
            in1 => \N__6512\,
            in2 => \N__6587\,
            in3 => \N__6391\,
            lcout => \Lab_UT.secuu0.un153_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_6_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__6513\,
            in1 => \N__6530\,
            in2 => \N__6421\,
            in3 => \N__6482\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13416\,
            ce => \N__6373\,
            sr => \N__12310\
        );

    \Lab_UT.secuu0.l_count_7_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__6483\,
            in1 => \N__6434\,
            in2 => \N__6395\,
            in3 => \N__6416\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13416\,
            ce => \N__6373\,
            sr => \N__12310\
        );

    \resetGen.reset_count_2_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100001"
        )
    port map (
            in0 => \N__6809\,
            in1 => \N__6719\,
            in2 => \N__6776\,
            in3 => \N__6753\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000001"
        )
    port map (
            in0 => \N__6754\,
            in1 => \N__6739\,
            in2 => \N__6727\,
            in3 => \N__6761\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__6802\,
            in1 => \N__6717\,
            in2 => \_gnd_net_\,
            in3 => \N__6752\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.un3_reset_count_i_a3_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__13463\,
            in1 => \N__10724\,
            in2 => \N__12172\,
            in3 => \N__7565\,
            lcout => \resetGen.N_104\,
            ltout => \resetGen.N_104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100000010"
        )
    port map (
            in0 => \N__6803\,
            in1 => \N__6718\,
            in2 => \N__6812\,
            in3 => \N__6788\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNO_0_2_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6787\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6800\,
            lcout => \resetGen.N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNITEEC1_2_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__6801\,
            in1 => \N__6786\,
            in2 => \_gnd_net_\,
            in3 => \N__6772\,
            lcout => \resetGen.N_86\,
            ltout => \resetGen.N_86_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000100"
        )
    port map (
            in0 => \N__6755\,
            in1 => \N__6740\,
            in2 => \N__6731\,
            in3 => \N__6723\,
            lcout => \resetGen.reset_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13411\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_44_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__11864\,
            in1 => \N__9704\,
            in2 => \N__9871\,
            in3 => \N__9965\,
            lcout => OPEN,
            ltout => \uu2.mem0.g2_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_25_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6845\,
            in2 => \N__6869\,
            in3 => \N__9440\,
            lcout => \uu2.mem0.g0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_40_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__9861\,
            in1 => \N__8473\,
            in2 => \_gnd_net_\,
            in3 => \N__8548\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_i_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_24_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__7688\,
            in1 => \N__11865\,
            in2 => \N__6860\,
            in3 => \N__12682\,
            lcout => \uu2.mem0.w_data_displaying_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_52_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9598\,
            in1 => \N__9540\,
            in2 => \N__9242\,
            in3 => \N__9162\,
            lcout => \uu2.mem0.g1_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_42_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000100101"
        )
    port map (
            in0 => \N__8547\,
            in1 => \N__12681\,
            in2 => \N__8477\,
            in3 => \N__12073\,
            lcout => \uu2.mem0.N_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_48_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011110"
        )
    port map (
            in0 => \N__12072\,
            in1 => \N__9869\,
            in2 => \N__12698\,
            in3 => \N__8417\,
            lcout => \uu2.mem0.g1_1_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_32_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111100011"
        )
    port map (
            in0 => \N__10936\,
            in1 => \N__10697\,
            in2 => \N__10625\,
            in3 => \N__11416\,
            lcout => \uu2.mem0.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_27_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000011"
        )
    port map (
            in0 => \N__8492\,
            in1 => \N__9705\,
            in2 => \N__6830\,
            in3 => \N__9964\,
            lcout => \uu2.mem0.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_60_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000110101011"
        )
    port map (
            in0 => \N__12370\,
            in1 => \N__9074\,
            in2 => \N__9257\,
            in3 => \N__9235\,
            lcout => \uu2.mem0.g0_i_6_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_38_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001111111"
        )
    port map (
            in0 => \N__9236\,
            in1 => \N__9062\,
            in2 => \N__7766\,
            in3 => \N__9164\,
            lcout => \uu2.mem0.g0_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_59_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__9800\,
            in1 => \N__9605\,
            in2 => \N__12371\,
            in3 => \N__9545\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_39_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__6899\,
            in1 => \N__8328\,
            in2 => \N__6893\,
            in3 => \N__9163\,
            lcout => \uu2.mem0.g0_i_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_53_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__11683\,
            in1 => \N__9422\,
            in2 => \N__9968\,
            in3 => \N__8546\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dicfsm.cState_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT_dicRun\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6944\,
            in2 => \N__6926\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7160\,
            in3 => \N__6878\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7443\,
            in1 => \N__6992\,
            in2 => \_gnd_net_\,
            in3 => \N__6875\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__13394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6976\,
            in2 => \_gnd_net_\,
            in3 => \N__6872\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__7445\,
            in1 => \N__7295\,
            in2 => \N__6962\,
            in3 => \N__7031\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNII0231_0_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__11794\,
            in1 => \N__7442\,
            in2 => \N__7300\,
            in3 => \N__7537\,
            lcout => \buart.Z_rx.bitcounte_0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__7444\,
            in1 => \N__7028\,
            in2 => \N__6980\,
            in3 => \N__7296\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_37_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__12694\,
            in1 => \N__8407\,
            in2 => \N__11244\,
            in3 => \N__8324\,
            lcout => \uu2.mem0.g0_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__7454\,
            in1 => \N__6924\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_RNIVHME_0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7858\,
            in1 => \N__7003\,
            in2 => \_gnd_net_\,
            in3 => \N__7538\,
            lcout => \buart.Z_rx.startbit\,
            ltout => \buart.Z_rx.startbit_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__6943\,
            in1 => \_gnd_net_\,
            in2 => \N__7007\,
            in3 => \N__6925\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_1_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7004\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6991\,
            in1 => \N__6975\,
            in2 => \N__6961\,
            in3 => \N__6942\,
            lcout => OPEN,
            ltout => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7155\,
            in2 => \N__6929\,
            in3 => \N__6923\,
            lcout => \buart.Z_rx.ser_clk\,
            ltout => \buart.Z_rx.ser_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__7156\,
            in1 => \N__7453\,
            in2 => \N__7169\,
            in3 => \N__7166\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_esr_0_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7142\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13385\,
            ce => \N__7253\,
            sr => \N__12302\
        );

    \uu2.r_data_reg_esr_1_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7127\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13385\,
            ce => \N__7253\,
            sr => \N__12302\
        );

    \uu2.r_data_reg_esr_2_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7112\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13385\,
            ce => \N__7253\,
            sr => \N__12302\
        );

    \uu2.r_data_reg_esr_3_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7097\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13385\,
            ce => \N__7253\,
            sr => \N__12302\
        );

    \uu2.r_data_reg_esr_4_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7085\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13385\,
            ce => \N__7253\,
            sr => \N__12302\
        );

    \uu2.r_data_reg_esr_5_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7073\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13385\,
            ce => \N__7253\,
            sr => \N__12302\
        );

    \uu2.r_data_reg_esr_6_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7049\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13385\,
            ce => \N__7253\,
            sr => \N__12302\
        );

    \uu2.r_data_reg_esr_7_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7274\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13385\,
            ce => \N__7253\,
            sr => \N__12302\
        );

    \buart.Z_tx.shifter_4_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__10277\,
            in1 => \N__7235\,
            in2 => \N__7217\,
            in3 => \N__10488\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13381\,
            ce => \N__8584\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_5_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__7229\,
            in1 => \N__10485\,
            in2 => \N__10289\,
            in3 => \N__7223\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13381\,
            ce => \N__8584\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_3_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__10276\,
            in1 => \N__7208\,
            in2 => \N__7202\,
            in3 => \N__10487\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13381\,
            ce => \N__8584\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_0_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__7841\,
            in1 => \N__10484\,
            in2 => \_gnd_net_\,
            in3 => \N__10278\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13381\,
            ce => \N__8584\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.uart_tx_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__10275\,
            in1 => \N__7193\,
            in2 => \_gnd_net_\,
            in3 => \N__10486\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13381\,
            ce => \N__8584\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10754\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7417\,
            in2 => \_gnd_net_\,
            in3 => \N__7172\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10821\,
            in2 => \_gnd_net_\,
            in3 => \N__7346\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10867\,
            in2 => \_gnd_net_\,
            in3 => \N__7343\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_4_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101101001110"
        )
    port map (
            in0 => \N__7517\,
            in1 => \N__7557\,
            in2 => \N__7478\,
            in3 => \N__7340\,
            lcout => \buart.Z_rx.bitcountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13414\,
            ce => \N__7391\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_0_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001011011110"
        )
    port map (
            in0 => \N__10761\,
            in1 => \N__7511\,
            in2 => \N__8892\,
            in3 => \N__7469\,
            lcout => \buart__rx_bitcount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13409\,
            ce => \N__7390\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_3_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100111100"
        )
    port map (
            in0 => \N__7468\,
            in1 => \N__10868\,
            in2 => \N__7337\,
            in3 => \N__7513\,
            lcout => \buart__rx_bitcount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13409\,
            ce => \N__7390\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_2_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001011011110"
        )
    port map (
            in0 => \N__10825\,
            in1 => \N__7512\,
            in2 => \N__7325\,
            in3 => \N__7470\,
            lcout => \buart__rx_bitcount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13409\,
            ce => \N__7390\,
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_15_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9035\,
            in1 => \N__11242\,
            in2 => \_gnd_net_\,
            in3 => \N__11984\,
            lcout => \uu2.mem0.w_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNI2B26_4_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10863\,
            in1 => \N__7559\,
            in2 => \N__7418\,
            in3 => \N__10819\,
            lcout => OPEN,
            ltout => \buart.Z_rx.N_103_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNIBJOC_0_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7304\,
            in2 => \N__7277\,
            in3 => \N__10753\,
            lcout => \buart.Z_rx.N_57_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNI8RI7_0_0_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10783\,
            in1 => \N__10760\,
            in2 => \N__10872\,
            in3 => \N__10818\,
            lcout => bu_rx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.un3_reset_count_i_a3_7_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__10820\,
            in1 => \N__12218\,
            in2 => \N__10873\,
            in3 => \N__10782\,
            lcout => \resetGen.un3_reset_count_i_a3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNIH513_4_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7558\,
            in2 => \_gnd_net_\,
            in3 => \N__7409\,
            lcout => \N_87\,
            ltout => \N_87_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNI8RI7_0_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__10817\,
            in1 => \N__10859\,
            in2 => \N__7541\,
            in3 => \N__10752\,
            lcout => \buart.Z_rx.N_91\,
            ltout => \buart.Z_rx.N_91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNIGM5F_0_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7520\,
            in3 => \N__11781\,
            lcout => \buart.Z_rx.N_29_0_i_2\,
            ltout => \buart.Z_rx.N_29_0_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_1_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011011110110"
        )
    port map (
            in0 => \N__7410\,
            in1 => \N__7493\,
            in2 => \N__7481\,
            in3 => \N__7474\,
            lcout => \buart.Z_rx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13403\,
            ce => \N__7383\,
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIAPHB1_5_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11848\,
            in1 => \N__12683\,
            in2 => \N__9872\,
            in3 => \N__12059\,
            lcout => \uu2.Z_decfrac105_7_3\,
            ltout => \uu2.Z_decfrac105_7_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011101100"
        )
    port map (
            in0 => \N__9371\,
            in1 => \N__11220\,
            in2 => \N__7358\,
            in3 => \N__10712\,
            lcout => \uu2.mem0.w_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_17_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7657\,
            in2 => \_gnd_net_\,
            in3 => \N__9369\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__11219\,
            in1 => \N__7706\,
            in2 => \N__7670\,
            in3 => \N__8230\,
            lcout => \uu2.mem0.w_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_18_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__12586\,
            in1 => \N__7658\,
            in2 => \_gnd_net_\,
            in3 => \N__9370\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011000"
        )
    port map (
            in0 => \N__11218\,
            in1 => \N__7697\,
            in2 => \N__7649\,
            in3 => \N__8231\,
            lcout => \uu2.mem0.w_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_5_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__12497\,
            in1 => \N__12792\,
            in2 => \N__11863\,
            in3 => \N__12685\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_5C_net\,
            ce => 'H',
            sr => \N__12281\
        );

    \uu2.w_addr_displaying_4_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__12684\,
            in1 => \N__12791\,
            in2 => \_gnd_net_\,
            in3 => \N__12498\,
            lcout => \uu2.w_addr_displayingZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_5C_net\,
            ce => 'H',
            sr => \N__12281\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__9280\,
            in1 => \N__11102\,
            in2 => \N__7622\,
            in3 => \N__11030\,
            lcout => \uu2.mem0.w_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_0_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8963\,
            in2 => \_gnd_net_\,
            in3 => \N__9320\,
            lcout => \uu2.un1_w_user_cr_0_0\,
            ltout => \uu2.un1_w_user_cr_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_wr_en_0_i_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110111011101"
        )
    port map (
            in0 => \N__7609\,
            in1 => \N__9279\,
            in2 => \N__7595\,
            in3 => \N__11101\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.rdy_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10154\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_34_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8180\,
            in1 => \N__8207\,
            in2 => \N__7745\,
            in3 => \N__7772\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_20_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9083\,
            in2 => \N__7730\,
            in3 => \N__7712\,
            lcout => OPEN,
            ltout => \uu2.mem0.un1_segment3_m6_0_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001100110"
        )
    port map (
            in0 => \N__11243\,
            in1 => \N__8216\,
            in2 => \N__7727\,
            in3 => \N__7676\,
            lcout => \uu2.mem0.w_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_35_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__8206\,
            in1 => \N__8179\,
            in2 => \_gnd_net_\,
            in3 => \N__7741\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_21_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001001000100"
        )
    port map (
            in0 => \N__10695\,
            in1 => \N__10617\,
            in2 => \N__11945\,
            in3 => \N__10943\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_22_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011001010"
        )
    port map (
            in0 => \N__10942\,
            in1 => \N__10696\,
            in2 => \N__10624\,
            in3 => \N__11462\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_rep1_RNI56RN_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__9410\,
            in1 => \N__8311\,
            in2 => \_gnd_net_\,
            in3 => \N__8520\,
            lcout => \uu2.g0_1_a5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_41_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8312\,
            in1 => \N__11564\,
            in2 => \N__12078\,
            in3 => \N__8406\,
            lcout => \uu2.mem0.g0_i_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_16_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__7757\,
            in1 => \N__9467\,
            in2 => \N__8264\,
            in3 => \N__8339\,
            lcout => \uu2.mem0.N_8_tz_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.g0_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13140\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13160\,
            lcout => OPEN,
            ltout => \led_c_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_56_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__9980\,
            in1 => \N__9699\,
            in2 => \N__7775\,
            in3 => \N__8429\,
            lcout => \uu2.mem0.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_58_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101000000"
        )
    port map (
            in0 => \N__9419\,
            in1 => \N__13161\,
            in2 => \N__13145\,
            in3 => \N__9148\,
            lcout => \uu2.mem0.g0_i_5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_30_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000010010"
        )
    port map (
            in0 => \N__8397\,
            in1 => \N__12693\,
            in2 => \N__9703\,
            in3 => \N__12065\,
            lcout => \uu2.mem0.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_rep1_8_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12798\,
            in1 => \N__9688\,
            in2 => \N__9763\,
            in3 => \N__8398\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_4_rep1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_8_rep1_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__12500\,
            in1 => \_gnd_net_\,
            in2 => \N__7751\,
            in3 => \N__8408\,
            lcout => \uu2.w_addr_displaying_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8_rep1C_net\,
            ce => 'H',
            sr => \N__12285\
        );

    \uu2.w_addr_displaying_8_rep1_RNIN6OC_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8309\,
            in2 => \_gnd_net_\,
            in3 => \N__8396\,
            lcout => OPEN,
            ltout => \uu2.N_42_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI8V6F2_3_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8594\,
            in1 => \N__12692\,
            in2 => \N__7748\,
            in3 => \N__12064\,
            lcout => \uu2.N_1482_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_7_rep1_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12802\,
            in1 => \N__12499\,
            in2 => \N__9764\,
            in3 => \N__8310\,
            lcout => \uu2.w_addr_displaying_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8_rep1C_net\,
            ce => 'H',
            sr => \N__12285\
        );

    \uu2.w_addr_displaying_4_rep1_RNI65VM_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__8308\,
            in1 => \N__9132\,
            in2 => \N__8409\,
            in3 => \N__9204\,
            lcout => \uu2.g0_1_a5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep1_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__9205\,
            in1 => \_gnd_net_\,
            in2 => \N__12808\,
            in3 => \N__12501\,
            lcout => \uu2.w_addr_displaying_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8_rep1C_net\,
            ce => 'H',
            sr => \N__12285\
        );

    \buart.Z_rx.shifter_7_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7859\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13380\,
            ce => \N__13255\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__7847\,
            in1 => \N__10517\,
            in2 => \N__7820\,
            in3 => \N__10279\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13378\,
            ce => \N__8583\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_2_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__7835\,
            in1 => \N__10518\,
            in2 => \N__7829\,
            in3 => \N__10280\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13378\,
            ce => \N__8583\,
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_4__un415_ci_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7927\,
            in1 => \N__8110\,
            in2 => \N__7803\,
            in3 => \N__11277\,
            lcout => \uu2.un415_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_2_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11280\,
            in1 => \N__7930\,
            in2 => \N__8119\,
            in3 => \N__8847\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__8777\
        );

    \uu2.vbuf_w_addr_user.result_1_3_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__7928\,
            in1 => \N__8111\,
            in2 => \N__7804\,
            in3 => \N__11278\,
            lcout => OPEN,
            ltout => \uu2.o_adder_vbuf_w_addr_user_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_3_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7799\,
            in2 => \N__7811\,
            in3 => \N__8846\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__8777\
        );

    \uu2.w_addr_user_RNIDD1A_5_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7792\,
            in1 => \N__7923\,
            in2 => \N__8032\,
            in3 => \N__11276\,
            lcout => \uu2.un2_w_addr_user_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_userZ0Z_1_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11279\,
            in1 => \N__7929\,
            in2 => \_gnd_net_\,
            in3 => \N__8845\,
            lcout => \uu2.w_addr_userZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_2C_net\,
            ce => 'H',
            sr => \N__8777\
        );

    \uu2.vbuf_w_addr_user.result_1_7_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__8140\,
            in1 => \N__7876\,
            in2 => \N__8085\,
            in3 => \N__7985\,
            lcout => OPEN,
            ltout => \uu2.o_adder_vbuf_w_addr_user_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_7_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8141\,
            in2 => \N__7901\,
            in3 => \N__8842\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_7C_net\,
            ce => 'H',
            sr => \N__8786\
        );

    \uu2.w_addr_user_6_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__8844\,
            in1 => \N__7877\,
            in2 => \N__8086\,
            in3 => \N__7987\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_7C_net\,
            ce => 'H',
            sr => \N__8786\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8138\,
            in1 => \N__11217\,
            in2 => \_gnd_net_\,
            in3 => \N__9706\,
            lcout => \uu2.mem0.w_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_8__un459_ci_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8074\,
            in2 => \_gnd_net_\,
            in3 => \N__8139\,
            lcout => OPEN,
            ltout => \uu2.vbuf_w_addr_user.un459_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.result_1_8_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__7875\,
            in1 => \N__7986\,
            in2 => \N__7883\,
            in3 => \N__8165\,
            lcout => OPEN,
            ltout => \uu2.o_adder_vbuf_w_addr_user_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_8_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__8166\,
            in1 => \_gnd_net_\,
            in2 => \N__7880\,
            in3 => \N__8843\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_7C_net\,
            ce => 'H',
            sr => \N__8786\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_6__un437_ci_3_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7968\,
            in2 => \_gnd_net_\,
            in3 => \N__8021\,
            lcout => \uu2.un437_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIKCH7_8_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__8167\,
            in1 => \N__8137\,
            in2 => \_gnd_net_\,
            in3 => \N__8115\,
            lcout => OPEN,
            ltout => \uu2.un2_w_addr_user_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIDMJM_4_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8081\,
            in1 => \N__7966\,
            in2 => \N__8048\,
            in3 => \N__8045\,
            lcout => \uu2.un2_w_addr_user\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.counter_gen_label_7__un448_ci_5_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9237\,
            in1 => \N__9582\,
            in2 => \_gnd_net_\,
            in3 => \N__9527\,
            lcout => \uu2.un448_ci_5\,
            ltout => \uu2.un448_ci_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_8_rep1_RNI5LHP1_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9463\,
            in1 => \N__8416\,
            in2 => \N__8036\,
            in3 => \N__8332\,
            lcout => \uu2.Z_decfrac106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_5_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__8855\,
            in1 => \N__7997\,
            in2 => \N__8031\,
            in3 => \N__7970\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__8781\
        );

    \uu2.w_addr_user_4_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__7996\,
            in1 => \N__7969\,
            in2 => \_gnd_net_\,
            in3 => \N__8854\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__8781\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7967\,
            in1 => \N__11201\,
            in2 => \_gnd_net_\,
            in3 => \N__12686\,
            lcout => \uu2.mem0.w_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_64_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9523\,
            in2 => \_gnd_net_\,
            in3 => \N__9155\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_46_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__12676\,
            in1 => \N__9870\,
            in2 => \N__7937\,
            in3 => \N__9361\,
            lcout => OPEN,
            ltout => \uu2.mem0.w_data_ns_1_1_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_26_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000111"
        )
    port map (
            in0 => \N__8741\,
            in1 => \N__11183\,
            in2 => \N__8234\,
            in3 => \N__8229\,
            lcout => \uu2.mem0.w_data_ns_1_0_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_5_rep1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__12677\,
            in1 => \N__12759\,
            in2 => \N__9539\,
            in3 => \N__12467\,
            lcout => \uu2.w_addr_displaying_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_5_rep1C_net\,
            ce => 'H',
            sr => \N__12282\
        );

    \uu2.w_addr_displaying_6_rep1_RNI6D891_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111111111"
        )
    port map (
            in0 => \N__9581\,
            in1 => \N__9522\,
            in2 => \N__12705\,
            in3 => \N__12049\,
            lcout => OPEN,
            ltout => \uu2.g0_1_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIRTT92_8_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010111"
        )
    port map (
            in0 => \N__12675\,
            in1 => \N__9695\,
            in2 => \N__8210\,
            in3 => \N__9957\,
            lcout => \uu2.g0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11999\,
            in1 => \N__12465\,
            in2 => \_gnd_net_\,
            in3 => \N__12050\,
            lcout => \uu2.w_addr_displayingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_5_rep1C_net\,
            ce => 'H',
            sr => \N__12282\
        );

    \uu2.w_addr_displaying_6_rep1_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101111010101010"
        )
    port map (
            in0 => \N__9589\,
            in1 => \N__9901\,
            in2 => \N__11825\,
            in3 => \N__12468\,
            lcout => \uu2.w_addr_displaying_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_5_rep1C_net\,
            ce => 'H',
            sr => \N__12282\
        );

    \uu2.w_addr_displaying_RNI2AJ42_5_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__9843\,
            in1 => \N__11847\,
            in2 => \N__8198\,
            in3 => \N__8189\,
            lcout => \uu2.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_rep1_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12462\,
            in1 => \N__11677\,
            in2 => \N__12601\,
            in3 => \N__9420\,
            lcout => \uu2.w_addr_displaying_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__12284\
        );

    \uu2.w_addr_displaying_2_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11676\,
            in1 => \N__12591\,
            in2 => \N__11592\,
            in3 => \N__12464\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__12284\
        );

    \uu2.w_addr_displaying_RNIUCHB1_2_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11571\,
            in1 => \N__11674\,
            in2 => \N__12600\,
            in3 => \N__12063\,
            lcout => \uu2.un15_w_data_displaying_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__11675\,
            in1 => \N__12590\,
            in2 => \_gnd_net_\,
            in3 => \N__12463\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__12284\
        );

    \uu2.w_addr_displaying_6_rep1_RNIAP701_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__8313\,
            in1 => \N__8399\,
            in2 => \N__9544\,
            in3 => \N__9603\,
            lcout => \uu2.g1_0_1\,
            ltout => \uu2.g1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_50_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100110011001"
        )
    port map (
            in0 => \N__9210\,
            in1 => \N__9135\,
            in2 => \N__8351\,
            in3 => \N__8251\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_28_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__8252\,
            in1 => \N__8240\,
            in2 => \N__8348\,
            in3 => \N__8345\,
            lcout => \uu2.mem0.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_51_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100100001001"
        )
    port map (
            in0 => \N__9209\,
            in1 => \N__9134\,
            in2 => \N__9966\,
            in3 => \N__8250\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_29_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__8314\,
            in1 => \_gnd_net_\,
            in2 => \N__8267\,
            in3 => \N__9604\,
            lcout => \uu2.mem0.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI7RCN_4_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000010001"
        )
    port map (
            in0 => \N__8521\,
            in1 => \N__9133\,
            in2 => \N__10019\,
            in3 => \N__8461\,
            lcout => \uu2.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_49_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__8462\,
            in1 => \N__9534\,
            in2 => \N__9421\,
            in3 => \N__9602\,
            lcout => \uu2.mem0.g1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_rep1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__12493\,
            in1 => \_gnd_net_\,
            in2 => \N__8534\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displaying_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0_rep1C_net\,
            ce => 'H',
            sr => \N__12286\
        );

    \uu2.mem0.ram512X8_inst_RNO_47_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000010001"
        )
    port map (
            in0 => \N__9136\,
            in1 => \N__8466\,
            in2 => \N__9228\,
            in3 => \N__8525\,
            lcout => \uu2.mem0.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_rep1_3_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__11586\,
            in1 => \N__11692\,
            in2 => \N__12602\,
            in3 => \N__9137\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_4_rep1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_rep1_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__9138\,
            in1 => \_gnd_net_\,
            in2 => \N__8480\,
            in3 => \N__12502\,
            lcout => \uu2.w_addr_displaying_3_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__12288\
        );

    \uu2.w_addr_displaying_1_rep1_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101001101010"
        )
    port map (
            in0 => \N__8467\,
            in1 => \N__12599\,
            in2 => \N__12509\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displaying_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__12288\
        );

    \uu2.w_addr_displaying_fast_2_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11693\,
            in1 => \N__12504\,
            in2 => \N__8441\,
            in3 => \N__12598\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__12288\
        );

    \uu2.mem0.ram512X8_inst_RNO_66_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110101111"
        )
    port map (
            in0 => \N__11633\,
            in1 => \N__8423\,
            in2 => \N__10018\,
            in3 => \N__8437\,
            lcout => \uu2.mem0.un1_segment4_0_i_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_4_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__10014\,
            in1 => \N__12503\,
            in2 => \_gnd_net_\,
            in3 => \N__12803\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1C_net\,
            ce => 'H',
            sr => \N__12288\
        );

    \uu2.mem0.ram512X8_inst_RNO_71_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__13030\,
            in1 => \N__12860\,
            in2 => \N__12983\,
            in3 => \N__13209\,
            lcout => \uu2.mem0.un1_segment4_0_i_i_a5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_RNIUTLC1_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__13210\,
            in1 => \N__13032\,
            in2 => \N__12876\,
            in3 => \N__12966\,
            lcout => \Lab_UT.didpuu0.didpsones.q13_0\,
            ltout => \Lab_UT.didpuu0.didpsones.q13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_2_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__10124\,
            in1 => \N__11732\,
            in2 => \N__8597\,
            in3 => \N__10076\,
            lcout => \Lab_UT_di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.g0_3_0_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001111101"
        )
    port map (
            in0 => \N__13208\,
            in1 => \N__12962\,
            in2 => \N__12875\,
            in3 => \N__13031\,
            lcout => \uu2.g0_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__8639\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8659\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8638\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.un1_bitcount_cry_0_c_RNO_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10236\,
            in1 => \N__10372\,
            in2 => \_gnd_net_\,
            in3 => \N__10317\,
            lcout => \buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIV5CT5_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10318\,
            in1 => \N__10509\,
            in2 => \_gnd_net_\,
            in3 => \N__10237\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_1_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__10516\,
            in1 => \N__10239\,
            in2 => \_gnd_net_\,
            in3 => \N__10028\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_0_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001100101001100"
        )
    port map (
            in0 => \N__10238\,
            in1 => \N__10371\,
            in2 => \N__10519\,
            in3 => \N__10319\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13382\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8637\,
            in2 => \N__8660\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8618\,
            in3 => \N__8723\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__13379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10324\,
            in1 => \N__8669\,
            in2 => \_gnd_net_\,
            in3 => \N__8720\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__13379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8696\,
            in3 => \N__8717\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__13379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__10325\,
            in1 => \_gnd_net_\,
            in2 => \N__8708\,
            in3 => \N__8714\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__13379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__8683\,
            in1 => \N__10323\,
            in2 => \_gnd_net_\,
            in3 => \N__8711\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13379\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8704\,
            in1 => \N__8692\,
            in2 => \N__8684\,
            in3 => \N__8668\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8655\,
            in1 => \N__8636\,
            in2 => \N__8617\,
            in3 => \N__8603\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_0_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11284\,
            in2 => \_gnd_net_\,
            in3 => \N__8853\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_0C_net\,
            ce => 'H',
            sr => \N__8785\
        );

    \uu2.w_addr_user_2_1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001011"
        )
    port map (
            in0 => \N__11905\,
            in1 => \N__8942\,
            in2 => \N__10691\,
            in3 => \N__11982\,
            lcout => OPEN,
            ltout => \uu2.w_addr_user_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNILAII7_4_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101110"
        )
    port map (
            in0 => \N__8921\,
            in1 => \N__10065\,
            in2 => \N__8792\,
            in3 => \N__11095\,
            lcout => OPEN,
            ltout => \uu2.w_addr_userZ2Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIT1MGD_4_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__8750\,
            in1 => \N__8927\,
            in2 => \N__8789\,
            in3 => \N__8807\,
            lcout => \uu2.w_addr_user_RNIT1MGDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_1_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001010"
        )
    port map (
            in0 => \N__10673\,
            in1 => \N__11354\,
            in2 => \N__10619\,
            in3 => \N__10918\,
            lcout => \uu2.w_addr_user_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNI24622_0_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__10920\,
            in1 => \N__8729\,
            in2 => \_gnd_net_\,
            in3 => \N__10143\,
            lcout => \Lab_UT.dspStr.cnt11_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dek.det_N_5_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__11983\,
            in1 => \N__11356\,
            in2 => \N__11420\,
            in3 => \N__11387\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrluu0.dek.det_NZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dek.det_N_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__11906\,
            in1 => \N__8936\,
            in2 => \N__8744\,
            in3 => \N__11457\,
            lcout => \Lab_UT.dicSelectLEDdisp\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_45_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110101"
        )
    port map (
            in0 => \N__10674\,
            in1 => \N__11355\,
            in2 => \N__10620\,
            in3 => \N__10919\,
            lcout => \uu2.mem0.N_1476_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un27_m3_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100001010"
        )
    port map (
            in0 => \N__10665\,
            in1 => \N__11357\,
            in2 => \N__10613\,
            in3 => \N__10917\,
            lcout => \uu2.un27_N_6_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNI11B71_3_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__13121\,
            in1 => \N__10595\,
            in2 => \N__11756\,
            in3 => \N__10666\,
            lcout => \Lab_UT.dspStr.cnt11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_m5_i_a3_2_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11455\,
            in1 => \N__11386\,
            in2 => \_gnd_net_\,
            in3 => \N__9053\,
            lcout => \uu2.w_m5_i_a3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dek.det_N_4_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11330\,
            in1 => \N__10769\,
            in2 => \_gnd_net_\,
            in3 => \N__11944\,
            lcout => \Lab_UT.dictrluu0.dek.det_NZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_0_0_0_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__11456\,
            in1 => \N__10916\,
            in2 => \_gnd_net_\,
            in3 => \N__11329\,
            lcout => OPEN,
            ltout => \uu2.un1_w_user_lf_0_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10591\,
            in2 => \N__8930\,
            in3 => \N__10664\,
            lcout => \uu2.un1_w_user_lf_2\,
            ltout => \uu2.un1_w_user_lf_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNILDNK6_4_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__8917\,
            in1 => \N__8803\,
            in2 => \N__8903\,
            in3 => \N__8900\,
            lcout => OPEN,
            ltout => \uu2.w_addr_user_RNILDNK6Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIOM3NG_4_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8893\,
            in2 => \N__8858\,
            in3 => \N__9017\,
            lcout => \uu2.un27_w_addr_user_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_5_a0_5_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9052\,
            in1 => \N__8982\,
            in2 => \N__9008\,
            in3 => \N__11382\,
            lcout => OPEN,
            ltout => \uu2.un1_w_user_lf_5_a0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_5_a0_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11409\,
            in2 => \N__8810\,
            in3 => \N__11882\,
            lcout => \uu2.un1_w_user_lf_5_aZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_1_rep1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11054\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT_dspStr_cnt_1_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13418\,
            ce => 'H',
            sr => \N__12303\
        );

    \Lab_UT.dspStr.cnt_2_rep1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11513\,
            lcout => \Lab_UT_dspStr_cnt_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13418\,
            ce => 'H',
            sr => \N__12303\
        );

    \Lab_UT.dspStr.cnt_3_rep1_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11306\,
            lcout => \Lab_UT_dspStr_cnt_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13418\,
            ce => 'H',
            sr => \N__12303\
        );

    \Lab_UT.dspStr.cnt_3_rep1_RNIIV651_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111001100"
        )
    port map (
            in0 => \N__8981\,
            in1 => \N__8999\,
            in2 => \N__11323\,
            in3 => \N__9050\,
            lcout => \Lab_UT_L3_tx_data_0_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_3_rep1_RNI05SQ_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__9051\,
            in1 => \_gnd_net_\,
            in2 => \N__9007\,
            in3 => \N__8980\,
            lcout => \Lab_UT_dspStr_un36_dOut\,
            ltout => \Lab_UT_dspStr_un36_dOut_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__11967\,
            in1 => \N__10963\,
            in2 => \N__9023\,
            in3 => \N__11023\,
            lcout => \uu2.un1_w_user_crZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un4_w_user_data_rdy_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__9292\,
            in1 => \N__11088\,
            in2 => \N__8959\,
            in3 => \N__9313\,
            lcout => \uu2.un4_w_user_data_rdyZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un27_m3_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101110011"
        )
    port map (
            in0 => \N__11448\,
            in1 => \N__10925\,
            in2 => \N__10618\,
            in3 => \N__8983\,
            lcout => OPEN,
            ltout => \uu2.un27_N_6_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un27_w_addr_user_i_1_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__9290\,
            in1 => \N__11086\,
            in2 => \N__9020\,
            in3 => \N__9311\,
            lcout => \uu2.un27_w_addr_user_iZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_3_rep1_RNIEPV31_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010100010"
        )
    port map (
            in0 => \N__10935\,
            in1 => \N__9006\,
            in2 => \N__11458\,
            in3 => \N__8984\,
            lcout => \L3_tx_data_0\,
            ltout => \L3_tx_data_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIQKOV8_8_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010101"
        )
    port map (
            in0 => \N__9291\,
            in1 => \N__11087\,
            in2 => \N__9323\,
            in3 => \N__9899\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_RNIQKOV8Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIB9CMF_8_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110101"
        )
    port map (
            in0 => \N__9312\,
            in1 => \N__9902\,
            in2 => \N__9296\,
            in3 => \N__9293\,
            lcout => \uu2.un21_w_addr_displaying_i\,
            ltout => \uu2.un21_w_addr_displaying_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_6_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101111111100000"
        )
    port map (
            in0 => \N__11817\,
            in1 => \N__9900\,
            in2 => \N__9260\,
            in3 => \N__12098\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_6C_net\,
            ce => 'H',
            sr => \N__12283\
        );

    \uu2.mem0.ram512X8_inst_RNO_69_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__12871\,
            in1 => \N__13055\,
            in2 => \N__12998\,
            in3 => \N__13226\,
            lcout => \uu2.mem0.g0_i_a11_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_55_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000100000"
        )
    port map (
            in0 => \N__13228\,
            in1 => \N__12991\,
            in2 => \N__13066\,
            in3 => \N__12874\,
            lcout => OPEN,
            ltout => \uu2.mem0.g3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_33_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010100000000"
        )
    port map (
            in0 => \N__12086\,
            in1 => \N__9238\,
            in2 => \N__9167\,
            in3 => \N__9156\,
            lcout => \uu2.mem0.un1_segment4_0_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_70_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__13225\,
            in1 => \N__12984\,
            in2 => \N__13065\,
            in3 => \N__12872\,
            lcout => \uu2.mem0.g0_i_a11_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_68_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__12873\,
            in1 => \_gnd_net_\,
            in2 => \N__12999\,
            in3 => \N__13227\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_i_a11_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_57_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111111111"
        )
    port map (
            in0 => \N__9616\,
            in1 => \N__11522\,
            in2 => \N__9065\,
            in3 => \N__9796\,
            lcout => \uu2.mem0.g0_i_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9617\,
            in2 => \_gnd_net_\,
            in3 => \N__12466\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_0C_net\,
            ce => 'H',
            sr => \N__12287\
        );

    \uu2.w_addr_displaying_fast_RNI3A1N_0_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__9615\,
            in1 => \N__9409\,
            in2 => \N__11637\,
            in3 => \N__9338\,
            lcout => \uu2.Z_decfrac106_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_61_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000010100"
        )
    port map (
            in0 => \N__11627\,
            in1 => \N__9787\,
            in2 => \N__12357\,
            in3 => \N__10006\,
            lcout => \uu2.mem0.bitmap_pmux_1_1_i_a5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_63_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9597\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9538\,
            lcout => OPEN,
            ltout => \uu2.mem0.g1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_43_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__9428\,
            in1 => \N__9476\,
            in2 => \N__9470\,
            in3 => \N__9462\,
            lcout => \uu2.mem0.g0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_62_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000010100"
        )
    port map (
            in0 => \N__10005\,
            in1 => \N__9411\,
            in2 => \N__9344\,
            in3 => \N__11628\,
            lcout => \uu2.mem0.bitmap_pmux_1_1_i_a5_2_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIFM1N_1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9412\,
            in1 => \N__9788\,
            in2 => \N__12358\,
            in3 => \N__9342\,
            lcout => \uu2.Z_decfrac105_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101001101010"
        )
    port map (
            in0 => \N__9343\,
            in1 => \N__12563\,
            in2 => \N__12508\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_1C_net\,
            ce => 'H',
            sr => \N__12289\
        );

    \uu2.w_addr_displaying_fast_3_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__11531\,
            in1 => \_gnd_net_\,
            in2 => \N__11638\,
            in3 => \N__12489\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_1C_net\,
            ce => 'H',
            sr => \N__12289\
        );

    \uu2.mem0.ram512X8_inst_RNO_65_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__10007\,
            in1 => \N__11629\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.mem0.Z_decfrac105_7_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_8_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12773\,
            in1 => \N__9671\,
            in2 => \N__9761\,
            in3 => \N__9944\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_4_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_8_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__9945\,
            in1 => \_gnd_net_\,
            in2 => \N__9971\,
            in3 => \N__12486\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \uu2.w_addr_displaying_RNI4K2N2_8_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12769\,
            in1 => \N__9669\,
            in2 => \N__9760\,
            in3 => \N__9943\,
            lcout => \uu2.un15_w_data_displaying\,
            ltout => \uu2.un15_w_data_displaying_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_6_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111011011001100"
        )
    port map (
            in0 => \N__11818\,
            in1 => \N__9842\,
            in2 => \N__9875\,
            in3 => \N__12487\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \uu2.w_addr_displaying_7_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12485\,
            in1 => \N__9750\,
            in2 => \N__12797\,
            in3 => \N__9672\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \uu2.w_addr_displaying_fast_7_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__12787\,
            in1 => \N__9795\,
            in2 => \N__9762\,
            in3 => \N__12488\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8C_net\,
            ce => 'H',
            sr => \N__12290\
        );

    \uu2.vbuf_w_addr_displaying.result_1_fast_8_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__12355\,
            in1 => \N__9749\,
            in2 => \N__12796\,
            in3 => \N__9670\,
            lcout => \uu2.w_addr_displaying_4_fast_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_RNO_0_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13223\,
            in2 => \N__11729\,
            in3 => \N__11730\,
            lcout => \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \Lab_UT.didpuu0.didpsones.un1_q_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_RNO_0_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12867\,
            in2 => \_gnd_net_\,
            in3 => \N__10127\,
            lcout => \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \Lab_UT.didpuu0.didpsones.un1_q_cry_0\,
            carryout => \Lab_UT.didpuu0.didpsones.un1_q_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_RNO_0_2_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13040\,
            in2 => \_gnd_net_\,
            in3 => \N__10118\,
            lcout => \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \Lab_UT.didpuu0.didpsones.un1_q_cry_1\,
            carryout => \Lab_UT.didpuu0.didpsones.un1_q_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_RNO_0_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12979\,
            in2 => \_gnd_net_\,
            in3 => \N__10115\,
            lcout => OPEN,
            ltout => \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_3_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__10079\,
            in1 => \N__10095\,
            in2 => \N__10112\,
            in3 => \N__11731\,
            lcout => \Lab_UT_di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_0_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__10109\,
            in1 => \N__11719\,
            in2 => \N__10096\,
            in3 => \N__10077\,
            lcout => \Lab_UT_di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_2_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010101010"
        )
    port map (
            in0 => \N__10532\,
            in1 => \_gnd_net_\,
            in2 => \N__10284\,
            in3 => \N__10505\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_1_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__10103\,
            in1 => \N__11720\,
            in2 => \N__10097\,
            in3 => \N__10078\,
            lcout => \Lab_UT_di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.un1_bitcount_cry_0_c_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10034\,
            in2 => \N__10373\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \buart.Z_tx.un1_bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10331\,
            in2 => \N__10352\,
            in3 => \N__10022\,
            lcout => \buart.Z_tx.bitcount_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \buart.Z_tx.un1_bitcount_cry_0\,
            carryout => \buart.Z_tx.un1_bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10400\,
            in2 => \N__10394\,
            in3 => \N__10526\,
            lcout => \buart.Z_tx.bitcount_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.un1_bitcount_cry_1\,
            carryout => \buart.Z_tx.un1_bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_3_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001111101100"
        )
    port map (
            in0 => \N__10244\,
            in1 => \N__10178\,
            in2 => \N__10523\,
            in3 => \N__10403\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIM5O32_2_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \N__10393\,
            in1 => \N__10240\,
            in2 => \_gnd_net_\,
            in3 => \N__10321\,
            lcout => \buart.Z_tx.bitcount_RNIM5O32Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIQOQA1_3_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10389\,
            in1 => \N__10347\,
            in2 => \N__10193\,
            in3 => \N__10367\,
            lcout => \buart__tx_uart_busy_0\,
            ltout => \buart__tx_uart_busy_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIL4O32_1_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \N__10348\,
            in1 => \_gnd_net_\,
            in2 => \N__10334\,
            in3 => \N__10320\,
            lcout => \buart.Z_tx.bitcount_RNIL4O32Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100001010"
        )
    port map (
            in0 => \N__10322\,
            in1 => \_gnd_net_\,
            in2 => \N__10274\,
            in3 => \N__10192\,
            lcout => \buart.Z_tx.un1_bitcount_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.sec_clkD_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13117\,
            lcout => \Lab_UT.sec_clkD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10144\,
            in2 => \N__10172\,
            in3 => \N__10168\,
            lcout => \Lab_UT.dspStr.cntZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \Lab_UT.dspStr.un1_cnt_3_cry_0\,
            clk => \N__13431\,
            ce => 'H',
            sr => \N__12306\
        );

    \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87E_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10924\,
            in2 => \_gnd_net_\,
            in3 => \N__10952\,
            lcout => \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87EZ0\,
            ltout => OPEN,
            carryin => \Lab_UT.dspStr.un1_cnt_3_cry_0\,
            carryout => \Lab_UT.dspStr.un1_cnt_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8E_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10679\,
            in2 => \_gnd_net_\,
            in3 => \N__10949\,
            lcout => \Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8EZ0\,
            ltout => OPEN,
            carryin => \Lab_UT.dspStr.un1_cnt_3_cry_1\,
            carryout => \Lab_UT.dspStr.un1_cnt_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9E_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10579\,
            in2 => \_gnd_net_\,
            in3 => \N__10946\,
            lcout => \Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9EZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_1_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11046\,
            lcout => \Lab_UT_dspStr_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13431\,
            ce => 'H',
            sr => \N__12306\
        );

    \Lab_UT.Lab3U01.q_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10763\,
            in1 => \N__10874\,
            in2 => \N__10829\,
            in3 => \N__10790\,
            lcout => \Lab_UT.rx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13428\,
            ce => 'H',
            sr => \N__12305\
        );

    \resetGen.un3_reset_count_i_a3_4_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__13511\,
            in1 => \N__13486\,
            in2 => \_gnd_net_\,
            in3 => \N__10762\,
            lcout => \resetGen.un3_reset_count_i_a3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNIN6202_3_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__10578\,
            in1 => \N__10675\,
            in2 => \_gnd_net_\,
            in3 => \N__11114\,
            lcout => \Lab_UT_L3_tx_data_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_2_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11502\,
            lcout => \Lab_UT_dspStr_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13428\,
            ce => 'H',
            sr => \N__12305\
        );

    \Lab_UT.dspStr.cnt_3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11298\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT_dspStr_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13428\,
            ce => 'H',
            sr => \N__12305\
        );

    \Lab_UT.dspStr.cnt_fast_3_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11299\,
            lcout => \Lab_UT.dspStr.cnt_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13428\,
            ce => 'H',
            sr => \N__12305\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11285\,
            in1 => \N__12584\,
            in2 => \_gnd_net_\,
            in3 => \N__11213\,
            lcout => \uu2.mem0.w_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_fast_RNIU9551_1_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001001011111"
        )
    port map (
            in0 => \N__11008\,
            in1 => \N__11934\,
            in2 => \N__11489\,
            in3 => \N__10987\,
            lcout => OPEN,
            ltout => \Lab_UT_L3_tx_data_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_4_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11066\,
            in1 => \N__11060\,
            in2 => \N__11117\,
            in3 => \N__11113\,
            lcout => \uu2.un1_w_user_crZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_fast_RNIQ5551_1_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110101111"
        )
    port map (
            in0 => \N__11007\,
            in1 => \N__11408\,
            in2 => \N__11488\,
            in3 => \N__10986\,
            lcout => \Lab_UT_L3_tx_data_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_fast_RNIS7551_1_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110110011"
        )
    port map (
            in0 => \N__11343\,
            in1 => \N__11005\,
            in2 => \N__10988\,
            in3 => \N__11476\,
            lcout => \Lab_UT_L3_tx_data_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_fast_1_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11053\,
            lcout => \Lab_UT.dspStr.cnt_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13425\,
            ce => 'H',
            sr => \N__12304\
        );

    \Lab_UT.dspStr.cnt_fast_RNIR6551_1_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000101"
        )
    port map (
            in0 => \N__10984\,
            in1 => \N__11378\,
            in2 => \N__11012\,
            in3 => \N__11483\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_fast_RNIT8551_1_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001111011011"
        )
    port map (
            in0 => \N__11006\,
            in1 => \N__10985\,
            in2 => \N__11487\,
            in3 => \N__11898\,
            lcout => \Lab_UT_L3_tx_data_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_fast_2_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11509\,
            lcout => \Lab_UT.dspStr.cnt_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13425\,
            ce => 'H',
            sr => \N__12304\
        );

    \Lab_UT.Lab3U00.q_esr_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12206\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT_rx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => \N__11765\,
            sr => \N__12300\
        );

    \Lab_UT.Lab3U00.q_esr_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12191\,
            lcout => \Lab_UT_rx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => \N__11765\,
            sr => \N__12300\
        );

    \Lab_UT.Lab3U00.q_esr_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT_rx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => \N__11765\,
            sr => \N__12300\
        );

    \Lab_UT.Lab3U00.q_esr_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13487\,
            lcout => \Lab_UT_rx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => \N__11765\,
            sr => \N__12300\
        );

    \Lab_UT.Lab3U00.q_esr_4_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13510\,
            lcout => \Lab_UT_rx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => \N__11765\,
            sr => \N__12300\
        );

    \Lab_UT.Lab3U00.q_esr_5_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12116\,
            lcout => \Lab_UT_rx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => \N__11765\,
            sr => \N__12300\
        );

    \Lab_UT.Lab3U00.q_esr_6_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12137\,
            lcout => \Lab_UT_rx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => \N__11765\,
            sr => \N__12300\
        );

    \Lab_UT.Lab3U00.q_esr_7_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12173\,
            lcout => \Lab_UT_rx_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13419\,
            ce => \N__11765\,
            sr => \N__12300\
        );

    \uu2.mem0.ram512X8_inst_RNO_54_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12097\,
            in2 => \_gnd_net_\,
            in3 => \N__12613\,
            lcout => \uu2.mem0.N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__11590\,
            in1 => \N__11695\,
            in2 => \N__12585\,
            in3 => \N__12080\,
            lcout => \uu2.w_addr_displaying_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_5_a0_4_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11966\,
            in1 => \N__11924\,
            in2 => \_gnd_net_\,
            in3 => \N__11899\,
            lcout => \uu2.un1_w_user_lf_5_a0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.counter_gen_label_6__un437_ci_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12804\,
            in1 => \N__11873\,
            in2 => \_gnd_net_\,
            in3 => \N__12706\,
            lcout => \uu2.un437_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.Lab3U00.q_esr_ctle_7_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11795\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12323\,
            lcout => \Lab_UT.Lab3U00.bu_rx_data_rdy_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.clkSecStrb_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13136\,
            in1 => \N__11755\,
            in2 => \_gnd_net_\,
            in3 => \N__13168\,
            lcout => \Lab_UT.didpuu0.clkSecStrbZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_fast_3_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11696\,
            in1 => \N__12561\,
            in2 => \N__11639\,
            in3 => \N__11591\,
            lcout => \uu2.w_addr_displaying_4_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_67_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010101000"
        )
    port map (
            in0 => \N__13054\,
            in1 => \N__12881\,
            in2 => \N__13000\,
            in3 => \N__13232\,
            lcout => \uu2.mem0.g0_i_a11_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_5_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__12495\,
            in1 => \N__12614\,
            in2 => \N__12809\,
            in3 => \N__12710\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_5C_net\,
            ce => 'H',
            sr => \N__12291\
        );

    \uu2.w_addr_displaying_0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12562\,
            in2 => \_gnd_net_\,
            in3 => \N__12496\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_5C_net\,
            ce => 'H',
            sr => \N__12291\
        );

    \uu2.w_addr_displaying_fast_8_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12494\,
            in1 => \N__12377\,
            in2 => \_gnd_net_\,
            in3 => \N__12356\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_5C_net\,
            ce => 'H',
            sr => \N__12291\
        );

    \resetGen.un3_reset_count_i_a3_5_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__12111\,
            in1 => \N__12186\,
            in2 => \N__12136\,
            in3 => \N__12202\,
            lcout => \resetGen.un3_reset_count_i_a3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13402\,
            ce => \N__13259\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13452\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13402\,
            ce => \N__13259\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_5_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12132\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13402\,
            ce => \N__13259\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_6_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12168\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13402\,
            ce => \N__13259\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_4_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12112\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13402\,
            ce => \N__13259\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_3_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13506\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13402\,
            ce => \N__13259\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_2_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13479\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13402\,
            ce => \N__13259\,
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.L3_led_1_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__12919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13224\,
            lcout => led_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.o_oneSecPluse_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13169\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13144\,
            lcout => led_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.L3_led_1_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12914\,
            in2 => \_gnd_net_\,
            in3 => \N__13067\,
            lcout => led_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.L3_led_1_3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__12915\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13001\,
            lcout => led_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.L3_led_1_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__12923\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12880\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Feb 28 2020 19:07:29

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15235\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15095\ : std_logic;
signal \N__15092\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal clk_in_c : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \Lab_UT.secuu0.un131_ci_3_cascade_\ : std_logic;
signal \Lab_UT.secuu0.un142_ci_0\ : std_logic;
signal \Lab_UT.secuu0.un131_ci_3\ : std_logic;
signal \Lab_UT.secuu0.un87_ci\ : std_logic;
signal \Lab_UT.secuu0.un87_ci_cascade_\ : std_logic;
signal \Lab_UT_L3_tx_data_0_4_cascade_\ : std_logic;
signal \Lab_UT_dspStr_un29_dOut_0_cascade_\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \Lab_UT.dspStr.un1_cnt_3_cry_0\ : std_logic;
signal \Lab_UT.dspStr.un1_cnt_3_cry_1\ : std_logic;
signal \Lab_UT.dspStr.un1_cnt_3_cry_2\ : std_logic;
signal \uu2.un1_w_user_lfZ0Z_4\ : std_logic;
signal \L3_tx_data_0_cascade_\ : std_logic;
signal \uu2.un1_w_user_lf_0\ : std_logic;
signal \uu2.un1_w_user_lf_0_cascade_\ : std_logic;
signal \INVuu2.w_addr_user_4C_net\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \uu2.un447_ci_3_cascade_\ : std_logic;
signal \uu2.o_adder_vbuf_w_addr_user_7\ : std_logic;
signal \uu2.mem0.w_addr_6\ : std_logic;
signal \uu2.mem0.w_addr_7\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \uu2.un447_ci_3\ : std_logic;
signal \uu2.vbuf_w_addr_user.un469_ci_0_cascade_\ : std_logic;
signal \uu2.o_adder_vbuf_w_addr_user_8\ : std_logic;
signal \Lab_UT.secuu0.un230_ci_1\ : std_logic;
signal \Lab_UT.secuu0.un109_ci\ : std_logic;
signal \Lab_UT.secuu0.un197_ci_9_cascade_\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_14\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_15\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_4\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_5\ : std_logic;
signal \Lab_UT.secuu0.l_precountZ0Z_3\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_1\ : std_logic;
signal \Lab_UT.secuu0.l_precountZ0Z_1\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_2\ : std_logic;
signal \Lab_UT.secuu0.l_precountZ0Z_2\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_0\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_14_cascade_\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_0_8\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_12\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_13\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_18_cascade_\ : std_logic;
signal \Lab_UT.dspStr.cnt11_1_cascade_\ : std_logic;
signal \Lab_UT.dspStr.cnt11_0_i\ : std_logic;
signal \Lab_UT.secuu0.un11_l_count_i\ : std_logic;
signal \Lab_UT_dspStr_un29_dOut_0\ : std_logic;
signal \uu2.un27_w_addr_user_0\ : std_logic;
signal \Lab_UT.dspStr.cntZ0Z_0\ : std_logic;
signal \uu2.un1_w_user_lfZ0Z_1\ : std_logic;
signal \uu2.un1_w_user_lfZ0Z_3\ : std_logic;
signal \uu2.un1_w_user_cr_0_0\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_2\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_2_cascade_\ : std_logic;
signal \uu2.un19_w_addr_userZ0Z_0_cascade_\ : std_logic;
signal \L3_tx_data_7\ : std_logic;
signal \uu2.mem0.w_data_7\ : std_logic;
signal \uu2.un1_w_user_cr_5Z0Z_1\ : std_logic;
signal \Lab_UT_L3_tx_data_2_0_cascade_\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_5\ : std_logic;
signal \Lab_UT_L3_tx_data_0_6\ : std_logic;
signal \uu2.mem0.w_data_6\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \uu2.mem0.w_addr_8\ : std_logic;
signal \Lab_UT_L3_tx_data_2_0\ : std_logic;
signal \uu2.mem0.w_addr_1\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \uu2.mem0.w_data_2\ : std_logic;
signal \uu2.un2_w_addr_user_5_cascade_\ : std_logic;
signal \uu2.un2_w_addr_user_4\ : std_logic;
signal \uu2.un2_w_addr_user\ : std_logic;
signal \uu2.un27_w_addr_user_i\ : std_logic;
signal \INVuu2.w_addr_user_3C_net\ : std_logic;
signal \uu2.w_addr_user_RNIKHHELZ0Z_2\ : std_logic;
signal \uu2.o_adder_vbuf_w_addr_user_3\ : std_logic;
signal \uu2.w_addr_userZ0Z_1\ : std_logic;
signal \uu2.un425_ci\ : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_10\ : std_logic;
signal \Lab_UT.secuu0.un186_ci_0_cascade_\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_8\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_9\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_7\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_3\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_11\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_11_cascade_\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_6\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_16\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_17\ : std_logic;
signal \Lab_UT.secuu0.un241_ci_2\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_16\ : std_logic;
signal \Lab_UT.secuu0.un263_ci\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_18\ : std_logic;
signal \Lab_UT.secuu0.un197_ci_9\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_12\ : std_logic;
signal \Lab_UT.secuu0.un153_ci\ : std_logic;
signal \Lab_UT.secuu0.un208_ci_0\ : std_logic;
signal \Lab_UT.secuu0.l_countZ0Z_13\ : std_logic;
signal \Lab_UT.secuu0.un11_l_count_i_g\ : std_logic;
signal \Lab_UT.secuu0.l_precountZ0Z_0\ : std_logic;
signal \uu2.un425_ci_0_cascade_\ : std_logic;
signal \uu2.vbuf_raddr.un469_ci_0_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \uu2.vbuf_raddr.un447_ci_3\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.vbuf_raddr.un447_ci_3_cascade_\ : std_logic;
signal \uu2.un425_ci_0\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_21\ : std_logic;
signal \uu2.mem0.w_data_0\ : std_logic;
signal \uu2.mem0.w_data_ns_1_5\ : std_logic;
signal \uu2.mem0.w_data_5\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_17\ : std_logic;
signal \uu2.mem0.G_14_0_a6_0_cascade_\ : std_logic;
signal \uu2.mem0.N_7_0_cascade_\ : std_logic;
signal \uu2.mem0.w_data_1\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_22\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_\ : std_logic;
signal \uu2.mem0.w_data_4\ : std_logic;
signal \uu2.mem0.G_14_0_a6_0_0_1\ : std_logic;
signal \uu2.mem0.w_data_3\ : std_logic;
signal \uu2.N_326_0_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_1_1_a8_1_2_0\ : std_logic;
signal \uu2.N_326_0\ : std_logic;
signal \uu2.bitmap_pmux_1_1_a8_1_1_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_1_1_a8_0_1\ : std_logic;
signal \uu2.bitmap_pmux_1_1_1_tz\ : std_logic;
signal \uu2.bitmap_pmux_1_1_1_tz_cascade_\ : std_logic;
signal \L3_tx_data_3\ : std_logic;
signal \uu2.mem0.w_data_1_0_0_3\ : std_logic;
signal \latticehx1k_pll_inst_PLLOUTCORE_i\ : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.mem0.w_addr_0\ : std_logic;
signal \INVuu2.w_addr_displaying_1C_net\ : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \buart.Z_rx.N_144_cascade_\ : std_logic;
signal \buart__rx_bitcount_4\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart__rx_bitcount_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \resetGen.reset_count_2_i_0_a3_5Z0Z_4_cascade_\ : std_logic;
signal bu_rx_data_5 : std_logic;
signal \resetGen.reset_count_2_i_0_a3_6Z0Z_4\ : std_logic;
signal \resetGen.reset_count_2_i_0_a3_4Z0Z_4\ : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal \buart.Z_rx.N_129_cascade_\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \buart.Z_rx.N_39\ : std_logic;
signal \Lab_UT_rx_data_4\ : std_logic;
signal \Lab_UT_rx_data_3\ : std_logic;
signal \Lab_UT.dictrluu0.N_103_1_cascade_\ : std_logic;
signal \Lab_UT_rx_data_5\ : std_logic;
signal \uu2.un1_w_user_lf_3Z0Z_1\ : std_logic;
signal \Lab_UT_dspStr_cnt_1\ : std_logic;
signal \Lab_UT_dspStr_cnt_3\ : std_logic;
signal \uu2.mem0.N_26_1_cascade_\ : std_logic;
signal \Lab_UT_dspStr_cnt_2\ : std_logic;
signal \Lab_UT.Lab3U00.bu_rx_data_rdy_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.mem0.w_addr_2\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.mem0.w_addr_3\ : std_logic;
signal \uu2.mem0.G_14_0_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_32_cascade_\ : std_logic;
signal \uu2.mem0.G_14_0_1\ : std_logic;
signal \uu2.N_329_0_cascade_\ : std_logic;
signal \uu2.Z_decfrac105_7\ : std_logic;
signal \N_52_0\ : std_logic;
signal \L3_segment2_0_0\ : std_logic;
signal \uu2.mem0.N_2159_0_cascade_\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_20\ : std_logic;
signal \L3_segment2_0\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4_cascade_\ : std_logic;
signal \uu2.mem0.g2_0\ : std_logic;
signal \uu2.mem0.N_5_cascade_\ : std_logic;
signal \uu2.mem0.bitmap_pmux_1_1_0_0\ : std_logic;
signal \uu2.mem0.N_14\ : std_logic;
signal \uu2.mem0.N_18\ : std_logic;
signal \uu2.mem0.un1_segment3_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_34\ : std_logic;
signal \uu2.Z_decfrac106\ : std_logic;
signal \uu2.mem0.un1_segment3_m2_1\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_47_cascade_\ : std_logic;
signal \uu2.mem0.un1_segment3_1_1\ : std_logic;
signal \uu2.mem0.N_2160_0\ : std_logic;
signal \N_52\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_48\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \uu2.mem0.w_addr_4\ : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \uu2.mem0.w_addr_5\ : std_logic;
signal \uu2.Z_decfrac106_2\ : std_logic;
signal \uu2.mem0.N_2160_1\ : std_logic;
signal \bfn_6_1_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.ser_clk_cascade_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal bu_rx_data_7 : std_logic;
signal bu_rx_data_6 : std_logic;
signal bu_rx_data_2 : std_logic;
signal bu_rx_data_4 : std_logic;
signal bu_rx_data_3 : std_logic;
signal \Lab_UT_rx_data_7\ : std_logic;
signal \Lab_UT_rx_data_1\ : std_logic;
signal \Lab_UT_rx_data_6\ : std_logic;
signal \Lab_UT.rx_data_rdy\ : std_logic;
signal \buart__rx_bitcount_0\ : std_logic;
signal \buart__rx_bitcount_2\ : std_logic;
signal \buart__rx_bitcount_3\ : std_logic;
signal \N_118\ : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \buart.Z_rx.ser_clk\ : std_logic;
signal \buart.Z_rx.N_129\ : std_logic;
signal \bu_rx_data_rdy_cascade_\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \buart.Z_rx.bitcount_e_0_RNII0231Z0Z_0\ : std_logic;
signal \Lab_UT_dec3_segmentUQ_0_6_cascade_\ : std_logic;
signal \N_71\ : std_logic;
signal \N_71_cascade_\ : std_logic;
signal \Lab_UT_dec3_segmentUQ_1_1_cascade_\ : std_logic;
signal \uu2.Z_decfrac105_7_2\ : std_logic;
signal \Lab_UT.rx_data_0\ : std_logic;
signal \Lab_UT.rx_dataZ0Z_2\ : std_logic;
signal \Lab_UT.dictrluu0.N_103_1\ : std_logic;
signal \Lab_UT.dicSelectLEDdisp\ : std_logic;
signal \Lab_UT.dicSelectLEDdisp_cascade_\ : std_logic;
signal \Lab_UT.dictrluu0.N_72\ : std_logic;
signal \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_o2_2\ : std_logic;
signal \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_3\ : std_logic;
signal \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_4\ : std_logic;
signal \Lab_UT.dictrluu0.dicfsm.N_102_cascade_\ : std_logic;
signal \uu2.N_93\ : std_logic;
signal \uu2.N_49_cascade_\ : std_logic;
signal \uu2.un1_segment3_m4_s_2\ : std_logic;
signal \uu2.g0_i_o4_0_1\ : std_logic;
signal \uu2.un1_segment3_m4_ns_1\ : std_logic;
signal \uu2.g0_i_o4_3_cascade_\ : std_logic;
signal \uu2.un1_segment3_m4\ : std_logic;
signal \uu2.w_addr_displaying_4_rep1_RNIMMRIAZ0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_53_cascade_\ : std_logic;
signal \uu2.mem0.un1_segment3_1_2\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4\ : std_logic;
signal \uu2.mem0.un1_segment3_m2_2\ : std_logic;
signal \uu2.mem0.un1_segment3_m2_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_42_cascade_\ : std_logic;
signal \uu2.mem0.un1_segment3_1_0\ : std_logic;
signal \Lab_UT.didpuu0.didpmtens.q_5_0_0_2\ : std_logic;
signal \uu2.un1_segment4_1_amZ0\ : std_logic;
signal \uu2.un1_segment4_1_bmZ0_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNIPN54Z0Z_8_cascade_\ : std_logic;
signal \uu2.N_292\ : std_logic;
signal \uu2.un1_segment4_5_amZ0Z_1\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNIV5694Z0Z_2\ : std_logic;
signal \uu2.N_290_0_i_0_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_RNI362A1Z0Z_3\ : std_logic;
signal \uu2.un1_w_addr_displaying_19_cascade_\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_\ : std_logic;
signal \uu2.mem0.N_5_0\ : std_logic;
signal \uu2.un1_segment3_s_0\ : std_logic;
signal \INVuu2.w_addr_displaying_5C_net\ : std_logic;
signal \uu2.un1_segment4_5_bmZ0\ : std_logic;
signal \Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMUZ0Z_0_cascade_\ : std_logic;
signal led_c_2 : std_logic;
signal \Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJZ0Z_0\ : std_logic;
signal \bfn_7_2_0_\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_0\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_1\ : std_logic;
signal \buart.Z_tx.un1_bitcount_axb_3\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_2\ : std_logic;
signal \buart.Z_tx.bitcount_RNIM5O32Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcount_RNIL4O32Z0Z_1\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \buart__tx_uart_busy_0_cascade_\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0\ : std_logic;
signal \resetGen.N_117\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \resetGen.N_117_cascade_\ : std_logic;
signal rst : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \resetGen.reset_countZ0Z_4\ : std_logic;
signal \resetGen.N_96_cascade_\ : std_logic;
signal \resetGen.N_133\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \buart__tx_uart_busy_0\ : std_logic;
signal \vbuf_tx_data_rdy_cascade_\ : std_logic;
signal \uu2.vbuf_tx_data_rdy_0\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal vbuf_tx_data_rdy : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \Lab_UT.secuu0.un4_l_count_0\ : std_logic;
signal \Lab_UT.secuu0.delay_lineZ0Z_0\ : std_logic;
signal \Lab_UT.secuu0.delay_lineZ0Z_1\ : std_logic;
signal \Lab_UT.didpuu0.didpmtens.N_122\ : std_logic;
signal \N_84_cascade_\ : std_logic;
signal \N_7\ : std_logic;
signal \uu2.un1_segment4_0_bmZ0\ : std_logic;
signal \uu2.un1_segment4_0_amZ0_cascade_\ : std_logic;
signal \uu2.un1_segment4_2_bmZ0\ : std_logic;
signal \uu2.un1_segment4_8_ns_1_cascade_\ : std_logic;
signal \uu2.un1_segment4_2_amZ0\ : std_logic;
signal \uu2.N_286\ : std_logic;
signal \Lab_UT.N_10_cascade_\ : std_logic;
signal \uu2.g0_i_o4_0_a8_2_2_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_5_rep1_RNIVO2EZ0Z1\ : std_logic;
signal \uu2.N_315_1_0\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_4C_net\ : std_logic;
signal \uu2.N_94\ : std_logic;
signal \uu2.bitmap_pmux_1_1_3_tz_1_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_1_1_3_tz\ : std_logic;
signal \uu2.N_111_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_4C_net\ : std_logic;
signal \uu2.un1_segment4_sn_N_36_mux_0_cascade_\ : std_logic;
signal \uu2.gZ0Z1\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_54\ : std_logic;
signal \uu2.un1_segment4_sn_N_58_0\ : std_logic;
signal \uu2.N_2150_0\ : std_logic;
signal \uu2.un1_segment4_sn_N_38_0_0\ : std_logic;
signal \uu2.g2_1_cascade_\ : std_logic;
signal \uu2.N_299_0\ : std_logic;
signal \uu2.un1_w_addr_displaying_inv_4_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_43\ : std_logic;
signal \uu2.segment3_m_1Z0Z_6_cascade_\ : std_logic;
signal \uu2.segment3_m_2_6_cascade_\ : std_logic;
signal \uu2.un1_segment4_4_bmZ0\ : std_logic;
signal \uu2.un1_segment4_4_amZ0_cascade_\ : std_logic;
signal \uu2.mem0.G_14_0_a6_2_1\ : std_logic;
signal \uu2.mem0.bitmap_pmux_1_1_2_tz_0\ : std_logic;
signal \uu2.bitmap_pmux_1_1_2_tz_1_0\ : std_logic;
signal \uu2.bitmap_pmux_1_1_2_tz_1_0_cascade_\ : std_logic;
signal \uu2.mem0.bitmap_pmux_1_1_2_tz_cascade_\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_33\ : std_logic;
signal \INVuu2.w_addr_displaying_2C_net\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \uu2.w_addr_displaying_RNI8NHB1Z0Z_2_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_RNI18582Z0Z_8\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.un3_r_clk_en_7\ : std_logic;
signal \uu2.un3_r_clk_en_0_0_cascade_\ : std_logic;
signal \uu2.un3_r_clk_en_6\ : std_logic;
signal \uu2_un3_r_clk_en_0_cascade_\ : std_logic;
signal \uu2.un349_ci_0\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.vbuf_count.un382_ci_8_1\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \uu2.un316_ci\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu2.un382_ci\ : std_logic;
signal uu2_un3_r_clk_en_0 : std_logic;
signal \uu2.l_countZ0Z_10\ : std_logic;
signal \Lab_UT.didpuu0.countEnMones_cascade_\ : std_logic;
signal \Lab_UT.didpuu0.didpmones.countEnMones_0\ : std_logic;
signal \Lab_UT.didpuu0.countEnStens_cascade_\ : std_logic;
signal \uu2.un1_segment4_2_amZ0Z_1\ : std_logic;
signal \uu2.w_addr_displaying_4_0_i_6_cascade_\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \uu2.g0_i_o4_0_a8_3_1\ : std_logic;
signal \uu2.w_addr_displaying_4_0_i_fast_6\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \uu2.un15_w_data_displaying_cascade_\ : std_logic;
signal \uu2.un19_w_addr_userZ0Z_0\ : std_logic;
signal \uu2.un21_w_addr_displaying_i_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_6C_net\ : std_logic;
signal \uu2.un15_w_data_displaying\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.w_addr_displaying_4_0_i_rep1_6\ : std_logic;
signal \uu2.w_addr_displaying_5_rep1_RNI3HMTZ0_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_6_rep1C_net\ : std_logic;
signal \uu2.un1_segment4_sn_N_61\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNI6N2KZ0Z_5_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNID5QHZ0Z_5\ : std_logic;
signal \uu2.un1_segment4_sn_N_39_0\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_RNILB202Z0Z_4\ : std_logic;
signal \uu2.N_92\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_3C_net\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNIN0TSZ0Z_4\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_4\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_2\ : std_logic;
signal \uu2.N_10_0\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.N_38\ : std_logic;
signal \Lab_UT.didpuu0.didpsones.N_32\ : std_logic;
signal \Lab_UT_dec0_un137_segmentUQ\ : std_logic;
signal \uu2.segment1_m_2Z0Z_0_cascade_\ : std_logic;
signal \uu2.segment1_m_0_cascade_\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_3\ : std_logic;
signal \uu2.segment3_m_6\ : std_logic;
signal \uu2.un1_segment1_iv_0_cascade_\ : std_logic;
signal \uu2.un1_segment1_0\ : std_logic;
signal \Lab_UT.didpuu0.didpstens.countEnStens_0\ : std_logic;
signal \uu2.un1_segment4_3_bmZ0\ : std_logic;
signal \uu2.un1_segment4_3_amZ0_cascade_\ : std_logic;
signal \uu2.un1_segment4_9_ns_1\ : std_logic;
signal \uu2.N_289_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNIFU9M8Z0Z_8\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_3\ : std_logic;
signal \uu2.N_1\ : std_logic;
signal \uu2.w_addr_displaying_4_rep1_RNIAVDBZ0Z_0\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNIKFIEZ0Z_6\ : std_logic;
signal \Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMUZ0Z_0_cascade_\ : std_logic;
signal led_c_3 : std_logic;
signal \Lab_UT.didpuu0.ledDisp00.selLed_RNI67CIZ0Z_0\ : std_logic;
signal \Lab_UT.un11_segmentUQ_1\ : std_logic;
signal \Lab_UT.didpuu0.countEnMtens_0_a4_0_cascade_\ : std_logic;
signal \Lab_UT.didpuu0.countEnMtens_0_a4_1\ : std_logic;
signal \Lab_UT.didpuu0.countEnMtens_0_a4_1_cascade_\ : std_logic;
signal \Lab_UT.didpuu0.countEnStens\ : std_logic;
signal \Lab_UT.didpuu0.countEnMtens\ : std_logic;
signal \Lab_UT.un152_segmentUQ_1\ : std_logic;
signal \Lab_UT.didpuu0.countEnMones\ : std_logic;
signal \uu2.un1_segment3_m5_bmZ0\ : std_logic;
signal bu_rx_data_1 : std_logic;
signal bu_rx_data_0 : std_logic;
signal \buart.Z_rx.N_41_i\ : std_logic;
signal clk_g : std_logic;
signal \Lab_UT.sec_clkD\ : std_logic;
signal \Lab_UT.didpuu0.clkSecStrbZ0\ : std_logic;
signal \L3_segment3_2\ : std_logic;
signal \L3_segment2_4_cascade_\ : std_logic;
signal \uu2.segment2_m_1Z0Z_6\ : std_logic;
signal \Lab_UT_di_Stens_2\ : std_logic;
signal \Lab_UT_di_Stens_3\ : std_logic;
signal \uu2.un1_segment3_m5_amZ0\ : std_logic;
signal \uu2.N_290_0_i_0\ : std_logic;
signal \uu2.un436_ci\ : std_logic;
signal \INVuu2.w_addr_displaying_4_rep1C_net\ : std_logic;
signal \uu2.w_addr_displaying_8_repZ0Z1\ : std_logic;
signal \uu2.un1_w_addr_displaying_35_0\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_4\ : std_logic;
signal \uu2.un1_w_addr_displaying_35_0_cascade_\ : std_logic;
signal \uu2.un1_w_addr_displaying_inv_2\ : std_logic;
signal \uu2.N_813_0_cascade_\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_58\ : std_logic;
signal \uu2.w_addr_displaying_7_repZ0Z1\ : std_logic;
signal \uu2.w_addr_displaying_4_repZ0Z1\ : std_logic;
signal \uu2.un1_segment3_m4_s_2_1\ : std_logic;
signal \Lab_UT_di_Sones_2\ : std_logic;
signal \Lab_UT_di_Sones_3\ : std_logic;
signal \uu2.un1_segment3_m0\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_6\ : std_logic;
signal \L3_segment1_3_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_5\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNIQD7R4Z0Z_5\ : std_logic;
signal \uu2.N_315_1\ : std_logic;
signal \uu2.w_addr_displaying_4_rep2_RNI75VMZ0\ : std_logic;
signal \uu2.un1_segment3_m5\ : std_logic;
signal \uu2.N_813_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_59\ : std_logic;
signal \uu2.segment2_m_2Z0Z_5\ : std_logic;
signal \uu2.segment2_m_5\ : std_logic;
signal \uu2.w_addr_displaying_0_repZ0Z1\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_7\ : std_logic;
signal \uu2.w_addr_displaying_4_rep2_RNI4S6JZ0\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNIEDBMZ0Z_7_cascade_\ : std_logic;
signal \uu2.un1_segment4_sn_N_38_0\ : std_logic;
signal \uu2.w_addr_displaying_4_repZ0Z2\ : std_logic;
signal \uu2.N_111\ : std_logic;
signal \uu2.w_addr_displaying_3_repZ0Z1\ : std_logic;
signal \uu2.Z_decfrac106_6\ : std_logic;
signal \uu2.un15_w_data_displaying_5\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_8\ : std_logic;
signal \INVuu2.w_addr_displaying_0_rep1C_net\ : std_logic;
signal \L3_segment4_2_cascade_\ : std_logic;
signal \uu2.N_280\ : std_logic;
signal \Lab_UT_di_Mtens_2\ : std_logic;
signal \Lab_UT_di_Mtens_3\ : std_logic;
signal \L3_segment4_4\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \INVuu2.w_addr_displaying_2_rep1C_net\ : std_logic;
signal \uu2.un1_w_addr_displaying_46_1\ : std_logic;
signal \uu2.un1_w_addr_displaying_46_1_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_RNI8U3D2Z0Z_0\ : std_logic;
signal \uu2.w_addr_displaying_5_repZ0Z1\ : std_logic;
signal \uu2.w_addr_displaying_6_repZ0Z1\ : std_logic;
signal \uu2.w_addr_displaying_2_repZ0Z1\ : std_logic;
signal \uu2.un1_w_addr_displaying_38_1\ : std_logic;
signal \uu2.segment3_m_3Z0Z_1\ : std_logic;
signal \uu2.un1_w_addr_displaying_38_1_cascade_\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \uu2.segment3_m_1\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.un21_w_addr_displaying_i\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_0\ : std_logic;
signal \INVuu2.w_addr_displaying_0C_net\ : std_logic;
signal rst_g : std_logic;
signal \uu2.mem0.N_2160_2\ : std_logic;
signal \Lab_UT_di_Sones_0\ : std_logic;
signal \Lab_UT_di_Stens_0\ : std_logic;
signal \Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11Z0Z_0_cascade_\ : std_logic;
signal led_c_0 : std_logic;
signal \Lab_UT_di_Mtens_0\ : std_logic;
signal \Lab_UT.didpuu0.ledDisp00.selLed_RNINURJZ0Z_0\ : std_logic;
signal \Lab_UT_di_Stens_1\ : std_logic;
signal \Lab_UT_di_Sones_1\ : std_logic;
signal \Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_1\ : std_logic;
signal led_c_1 : std_logic;
signal \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_0\ : std_logic;
signal \Lab_UT_di_Mtens_1\ : std_logic;
signal \Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJZ0Z_0\ : std_logic;
signal \Lab_UT_di_Mones_2\ : std_logic;
signal \Lab_UT_di_Mones_1\ : std_logic;
signal \Lab_UT_di_Mones_3\ : std_logic;
signal \Lab_UT_di_Mones_0\ : std_logic;
signal \uu2.N_2160_1_0_0\ : std_logic;
signal \Lab_UT_dicRun\ : std_logic;
signal \Lab_UT_l_oneSecPluse\ : std_logic;
signal led_c_4 : std_logic;
signal \_gnd_net_\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__7968\&\N__7830\&\N__7878\&\N__7950\&\N__7920\&\N__7806\&\N__11109\&\N__11322\&\N__11283\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__6996\&\N__6495\&\N__6510\&\N__9297\&\N__9342\&\N__8964\&\N__9009\&\N__6981\&\N__8058\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&\N__6870\&'0'&\N__7026\&'0'&\N__7752\&'0'&\N__7995\&'0'&\N__7980\&'0'&\N__6948\&'0'&\N__8013\&'0'&\N__7770\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \latticehx1k_pll_inst_PLLOUTCORE_i\,
            REFERENCECLK => \N__6339\,
            RESETB => \N__8370\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => \N__11235\,
            RCLK => \N__13508\,
            RE => \N__11232\,
            WCLKE => \N__8121\,
            WCLK => \N__13509\,
            WE => \N__8120\
        );

    \led_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17566\,
            DIN => \N__17565\,
            DOUT => \N__17564\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17566\,
            PADOUT => \N__17565\,
            PADIN => \N__17564\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16500\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17557\,
            DIN => \N__17556\,
            DOUT => \N__17555\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17557\,
            PADOUT => \N__17556\,
            PADIN => \N__17555\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17127\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17548\,
            DIN => \N__17547\,
            DOUT => \N__17546\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17548\,
            PADOUT => \N__17547\,
            PADIN => \N__17546\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8232\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17539\,
            DIN => \N__17538\,
            DOUT => \N__17537\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17539\,
            PADOUT => \N__17538\,
            PADIN => \N__17537\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17530\,
            DIN => \N__17529\,
            DOUT => \N__17528\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17530\,
            PADOUT => \N__17529\,
            PADIN => \N__17528\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10611\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17521\,
            DIN => \N__17520\,
            DOUT => \N__17519\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17521\,
            PADOUT => \N__17520\,
            PADIN => \N__17519\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13263\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17512\,
            DIN => \N__17511\,
            DOUT => \N__17510\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17512\,
            PADOUT => \N__17511\,
            PADIN => \N__17510\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17463\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17503\,
            DIN => \N__17502\,
            DOUT => \N__17501\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__17503\,
            PADOUT => \N__17502\,
            PADIN => \N__17501\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__13514\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17494\,
            DIN => \N__17493\,
            DOUT => \N__17492\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__17494\,
            PADOUT => \N__17493\,
            PADIN => \N__17492\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17485\,
            DIN => \N__17484\,
            DOUT => \N__17483\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17485\,
            PADOUT => \N__17484\,
            PADIN => \N__17483\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__4248\ : CascadeMux
    port map (
            O => \N__17466\,
            I => \Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11Z0Z_0_cascade_\
        );

    \I__4247\ : IoInMux
    port map (
            O => \N__17463\,
            I => \N__17460\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__17460\,
            I => \N__17457\
        );

    \I__4245\ : Span12Mux_s3_h
    port map (
            O => \N__17457\,
            I => \N__17454\
        );

    \I__4244\ : Odrv12
    port map (
            O => \N__17454\,
            I => led_c_0
        );

    \I__4243\ : InMux
    port map (
            O => \N__17451\,
            I => \N__17444\
        );

    \I__4242\ : InMux
    port map (
            O => \N__17450\,
            I => \N__17439\
        );

    \I__4241\ : InMux
    port map (
            O => \N__17449\,
            I => \N__17436\
        );

    \I__4240\ : InMux
    port map (
            O => \N__17448\,
            I => \N__17431\
        );

    \I__4239\ : InMux
    port map (
            O => \N__17447\,
            I => \N__17431\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__17444\,
            I => \N__17428\
        );

    \I__4237\ : InMux
    port map (
            O => \N__17443\,
            I => \N__17423\
        );

    \I__4236\ : InMux
    port map (
            O => \N__17442\,
            I => \N__17423\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__17439\,
            I => \N__17412\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__17436\,
            I => \N__17409\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__17431\,
            I => \N__17406\
        );

    \I__4232\ : Span4Mux_v
    port map (
            O => \N__17428\,
            I => \N__17401\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__17423\,
            I => \N__17401\
        );

    \I__4230\ : CascadeMux
    port map (
            O => \N__17422\,
            I => \N__17397\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__17421\,
            I => \N__17394\
        );

    \I__4228\ : InMux
    port map (
            O => \N__17420\,
            I => \N__17390\
        );

    \I__4227\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17379\
        );

    \I__4226\ : InMux
    port map (
            O => \N__17418\,
            I => \N__17379\
        );

    \I__4225\ : InMux
    port map (
            O => \N__17417\,
            I => \N__17379\
        );

    \I__4224\ : InMux
    port map (
            O => \N__17416\,
            I => \N__17379\
        );

    \I__4223\ : InMux
    port map (
            O => \N__17415\,
            I => \N__17379\
        );

    \I__4222\ : Span4Mux_h
    port map (
            O => \N__17412\,
            I => \N__17370\
        );

    \I__4221\ : Span4Mux_v
    port map (
            O => \N__17409\,
            I => \N__17370\
        );

    \I__4220\ : Span4Mux_v
    port map (
            O => \N__17406\,
            I => \N__17370\
        );

    \I__4219\ : Span4Mux_v
    port map (
            O => \N__17401\,
            I => \N__17370\
        );

    \I__4218\ : InMux
    port map (
            O => \N__17400\,
            I => \N__17363\
        );

    \I__4217\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17363\
        );

    \I__4216\ : InMux
    port map (
            O => \N__17394\,
            I => \N__17363\
        );

    \I__4215\ : InMux
    port map (
            O => \N__17393\,
            I => \N__17360\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__17390\,
            I => \Lab_UT_di_Mtens_0\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__17379\,
            I => \Lab_UT_di_Mtens_0\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__17370\,
            I => \Lab_UT_di_Mtens_0\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__17363\,
            I => \Lab_UT_di_Mtens_0\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__17360\,
            I => \Lab_UT_di_Mtens_0\
        );

    \I__4209\ : InMux
    port map (
            O => \N__17349\,
            I => \N__17346\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__17346\,
            I => \Lab_UT.didpuu0.ledDisp00.selLed_RNINURJZ0Z_0\
        );

    \I__4207\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17339\
        );

    \I__4206\ : InMux
    port map (
            O => \N__17342\,
            I => \N__17336\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__17339\,
            I => \N__17332\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__17336\,
            I => \N__17322\
        );

    \I__4203\ : InMux
    port map (
            O => \N__17335\,
            I => \N__17319\
        );

    \I__4202\ : Span4Mux_h
    port map (
            O => \N__17332\,
            I => \N__17313\
        );

    \I__4201\ : InMux
    port map (
            O => \N__17331\,
            I => \N__17310\
        );

    \I__4200\ : InMux
    port map (
            O => \N__17330\,
            I => \N__17303\
        );

    \I__4199\ : InMux
    port map (
            O => \N__17329\,
            I => \N__17303\
        );

    \I__4198\ : InMux
    port map (
            O => \N__17328\,
            I => \N__17303\
        );

    \I__4197\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17300\
        );

    \I__4196\ : InMux
    port map (
            O => \N__17326\,
            I => \N__17294\
        );

    \I__4195\ : InMux
    port map (
            O => \N__17325\,
            I => \N__17294\
        );

    \I__4194\ : Span4Mux_v
    port map (
            O => \N__17322\,
            I => \N__17289\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__17319\,
            I => \N__17289\
        );

    \I__4192\ : InMux
    port map (
            O => \N__17318\,
            I => \N__17284\
        );

    \I__4191\ : InMux
    port map (
            O => \N__17317\,
            I => \N__17284\
        );

    \I__4190\ : InMux
    port map (
            O => \N__17316\,
            I => \N__17281\
        );

    \I__4189\ : Sp12to4
    port map (
            O => \N__17313\,
            I => \N__17272\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__17310\,
            I => \N__17272\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__17303\,
            I => \N__17272\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__17300\,
            I => \N__17272\
        );

    \I__4185\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17269\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__17294\,
            I => \Lab_UT_di_Stens_1\
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__17289\,
            I => \Lab_UT_di_Stens_1\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__17284\,
            I => \Lab_UT_di_Stens_1\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__17281\,
            I => \Lab_UT_di_Stens_1\
        );

    \I__4180\ : Odrv12
    port map (
            O => \N__17272\,
            I => \Lab_UT_di_Stens_1\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__17269\,
            I => \Lab_UT_di_Stens_1\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__17256\,
            I => \N__17249\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__17255\,
            I => \N__17243\
        );

    \I__4176\ : InMux
    port map (
            O => \N__17254\,
            I => \N__17240\
        );

    \I__4175\ : InMux
    port map (
            O => \N__17253\,
            I => \N__17234\
        );

    \I__4174\ : InMux
    port map (
            O => \N__17252\,
            I => \N__17225\
        );

    \I__4173\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17225\
        );

    \I__4172\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17225\
        );

    \I__4171\ : InMux
    port map (
            O => \N__17247\,
            I => \N__17225\
        );

    \I__4170\ : InMux
    port map (
            O => \N__17246\,
            I => \N__17220\
        );

    \I__4169\ : InMux
    port map (
            O => \N__17243\,
            I => \N__17220\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__17240\,
            I => \N__17217\
        );

    \I__4167\ : InMux
    port map (
            O => \N__17239\,
            I => \N__17214\
        );

    \I__4166\ : CascadeMux
    port map (
            O => \N__17238\,
            I => \N__17211\
        );

    \I__4165\ : InMux
    port map (
            O => \N__17237\,
            I => \N__17206\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__17234\,
            I => \N__17201\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__17225\,
            I => \N__17201\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__17220\,
            I => \N__17198\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__17217\,
            I => \N__17193\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__17214\,
            I => \N__17193\
        );

    \I__4159\ : InMux
    port map (
            O => \N__17211\,
            I => \N__17186\
        );

    \I__4158\ : InMux
    port map (
            O => \N__17210\,
            I => \N__17186\
        );

    \I__4157\ : InMux
    port map (
            O => \N__17209\,
            I => \N__17186\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__17206\,
            I => \N__17183\
        );

    \I__4155\ : Span4Mux_v
    port map (
            O => \N__17201\,
            I => \N__17178\
        );

    \I__4154\ : Span4Mux_v
    port map (
            O => \N__17198\,
            I => \N__17178\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__17193\,
            I => \Lab_UT_di_Sones_1\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__17186\,
            I => \Lab_UT_di_Sones_1\
        );

    \I__4151\ : Odrv12
    port map (
            O => \N__17183\,
            I => \Lab_UT_di_Sones_1\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__17178\,
            I => \Lab_UT_di_Sones_1\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__17169\,
            I => \Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11Z0Z_0_cascade_\
        );

    \I__4148\ : InMux
    port map (
            O => \N__17166\,
            I => \N__17159\
        );

    \I__4147\ : InMux
    port map (
            O => \N__17165\,
            I => \N__17159\
        );

    \I__4146\ : InMux
    port map (
            O => \N__17164\,
            I => \N__17156\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__17159\,
            I => \N__17151\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__17156\,
            I => \N__17151\
        );

    \I__4143\ : Span4Mux_h
    port map (
            O => \N__17151\,
            I => \N__17147\
        );

    \I__4142\ : InMux
    port map (
            O => \N__17150\,
            I => \N__17144\
        );

    \I__4141\ : Span4Mux_v
    port map (
            O => \N__17147\,
            I => \N__17140\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__17144\,
            I => \N__17137\
        );

    \I__4139\ : InMux
    port map (
            O => \N__17143\,
            I => \N__17134\
        );

    \I__4138\ : Odrv4
    port map (
            O => \N__17140\,
            I => \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_1\
        );

    \I__4137\ : Odrv12
    port map (
            O => \N__17137\,
            I => \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_1\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__17134\,
            I => \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_1\
        );

    \I__4135\ : IoInMux
    port map (
            O => \N__17127\,
            I => \N__17124\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__17124\,
            I => \N__17121\
        );

    \I__4133\ : Span4Mux_s3_h
    port map (
            O => \N__17121\,
            I => \N__17118\
        );

    \I__4132\ : Odrv4
    port map (
            O => \N__17118\,
            I => led_c_1
        );

    \I__4131\ : InMux
    port map (
            O => \N__17115\,
            I => \N__17101\
        );

    \I__4130\ : InMux
    port map (
            O => \N__17114\,
            I => \N__17101\
        );

    \I__4129\ : InMux
    port map (
            O => \N__17113\,
            I => \N__17101\
        );

    \I__4128\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17101\
        );

    \I__4127\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17098\
        );

    \I__4126\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17095\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__17101\,
            I => \N__17086\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__17098\,
            I => \N__17086\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__17095\,
            I => \N__17086\
        );

    \I__4122\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17081\
        );

    \I__4121\ : InMux
    port map (
            O => \N__17093\,
            I => \N__17081\
        );

    \I__4120\ : Span12Mux_s6_h
    port map (
            O => \N__17086\,
            I => \N__17074\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__17081\,
            I => \N__17074\
        );

    \I__4118\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17069\
        );

    \I__4117\ : InMux
    port map (
            O => \N__17079\,
            I => \N__17069\
        );

    \I__4116\ : Odrv12
    port map (
            O => \N__17074\,
            I => \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_0\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__17069\,
            I => \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_0\
        );

    \I__4114\ : InMux
    port map (
            O => \N__17064\,
            I => \N__17058\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__17063\,
            I => \N__17055\
        );

    \I__4112\ : InMux
    port map (
            O => \N__17062\,
            I => \N__17051\
        );

    \I__4111\ : InMux
    port map (
            O => \N__17061\,
            I => \N__17046\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__17058\,
            I => \N__17040\
        );

    \I__4109\ : InMux
    port map (
            O => \N__17055\,
            I => \N__17035\
        );

    \I__4108\ : InMux
    port map (
            O => \N__17054\,
            I => \N__17035\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__17051\,
            I => \N__17032\
        );

    \I__4106\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17027\
        );

    \I__4105\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17027\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__17046\,
            I => \N__17024\
        );

    \I__4103\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17017\
        );

    \I__4102\ : InMux
    port map (
            O => \N__17044\,
            I => \N__17017\
        );

    \I__4101\ : InMux
    port map (
            O => \N__17043\,
            I => \N__17017\
        );

    \I__4100\ : Span4Mux_v
    port map (
            O => \N__17040\,
            I => \N__17014\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__17035\,
            I => \N__17011\
        );

    \I__4098\ : Span4Mux_v
    port map (
            O => \N__17032\,
            I => \N__17006\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__17027\,
            I => \N__17006\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__17024\,
            I => \N__16991\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__17017\,
            I => \N__16991\
        );

    \I__4094\ : Span4Mux_h
    port map (
            O => \N__17014\,
            I => \N__16991\
        );

    \I__4093\ : Span4Mux_v
    port map (
            O => \N__17011\,
            I => \N__16991\
        );

    \I__4092\ : Span4Mux_v
    port map (
            O => \N__17006\,
            I => \N__16991\
        );

    \I__4091\ : InMux
    port map (
            O => \N__17005\,
            I => \N__16982\
        );

    \I__4090\ : InMux
    port map (
            O => \N__17004\,
            I => \N__16982\
        );

    \I__4089\ : InMux
    port map (
            O => \N__17003\,
            I => \N__16982\
        );

    \I__4088\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16982\
        );

    \I__4087\ : Odrv4
    port map (
            O => \N__16991\,
            I => \Lab_UT_di_Mtens_1\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__16982\,
            I => \Lab_UT_di_Mtens_1\
        );

    \I__4085\ : InMux
    port map (
            O => \N__16977\,
            I => \N__16974\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__16974\,
            I => \Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJZ0Z_0\
        );

    \I__4083\ : InMux
    port map (
            O => \N__16971\,
            I => \N__16967\
        );

    \I__4082\ : InMux
    port map (
            O => \N__16970\,
            I => \N__16960\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__16967\,
            I => \N__16957\
        );

    \I__4080\ : InMux
    port map (
            O => \N__16966\,
            I => \N__16954\
        );

    \I__4079\ : CascadeMux
    port map (
            O => \N__16965\,
            I => \N__16950\
        );

    \I__4078\ : CascadeMux
    port map (
            O => \N__16964\,
            I => \N__16947\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__16963\,
            I => \N__16943\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__16960\,
            I => \N__16940\
        );

    \I__4075\ : Span4Mux_v
    port map (
            O => \N__16957\,
            I => \N__16933\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__16954\,
            I => \N__16933\
        );

    \I__4073\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16917\
        );

    \I__4072\ : InMux
    port map (
            O => \N__16950\,
            I => \N__16917\
        );

    \I__4071\ : InMux
    port map (
            O => \N__16947\,
            I => \N__16917\
        );

    \I__4070\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16917\
        );

    \I__4069\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16917\
        );

    \I__4068\ : Span4Mux_v
    port map (
            O => \N__16940\,
            I => \N__16914\
        );

    \I__4067\ : InMux
    port map (
            O => \N__16939\,
            I => \N__16911\
        );

    \I__4066\ : InMux
    port map (
            O => \N__16938\,
            I => \N__16908\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__16933\,
            I => \N__16905\
        );

    \I__4064\ : InMux
    port map (
            O => \N__16932\,
            I => \N__16902\
        );

    \I__4063\ : InMux
    port map (
            O => \N__16931\,
            I => \N__16893\
        );

    \I__4062\ : InMux
    port map (
            O => \N__16930\,
            I => \N__16893\
        );

    \I__4061\ : InMux
    port map (
            O => \N__16929\,
            I => \N__16893\
        );

    \I__4060\ : InMux
    port map (
            O => \N__16928\,
            I => \N__16893\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__16917\,
            I => \N__16890\
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__16914\,
            I => \Lab_UT_di_Mones_2\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__16911\,
            I => \Lab_UT_di_Mones_2\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__16908\,
            I => \Lab_UT_di_Mones_2\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__16905\,
            I => \Lab_UT_di_Mones_2\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__16902\,
            I => \Lab_UT_di_Mones_2\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__16893\,
            I => \Lab_UT_di_Mones_2\
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__16890\,
            I => \Lab_UT_di_Mones_2\
        );

    \I__4051\ : InMux
    port map (
            O => \N__16875\,
            I => \N__16870\
        );

    \I__4050\ : InMux
    port map (
            O => \N__16874\,
            I => \N__16867\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__16873\,
            I => \N__16856\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__16870\,
            I => \N__16852\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__16867\,
            I => \N__16849\
        );

    \I__4046\ : CascadeMux
    port map (
            O => \N__16866\,
            I => \N__16845\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__16865\,
            I => \N__16842\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__16864\,
            I => \N__16837\
        );

    \I__4043\ : InMux
    port map (
            O => \N__16863\,
            I => \N__16826\
        );

    \I__4042\ : InMux
    port map (
            O => \N__16862\,
            I => \N__16826\
        );

    \I__4041\ : InMux
    port map (
            O => \N__16861\,
            I => \N__16826\
        );

    \I__4040\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16826\
        );

    \I__4039\ : InMux
    port map (
            O => \N__16859\,
            I => \N__16826\
        );

    \I__4038\ : InMux
    port map (
            O => \N__16856\,
            I => \N__16821\
        );

    \I__4037\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16821\
        );

    \I__4036\ : Span4Mux_v
    port map (
            O => \N__16852\,
            I => \N__16816\
        );

    \I__4035\ : Span4Mux_v
    port map (
            O => \N__16849\,
            I => \N__16816\
        );

    \I__4034\ : InMux
    port map (
            O => \N__16848\,
            I => \N__16813\
        );

    \I__4033\ : InMux
    port map (
            O => \N__16845\,
            I => \N__16802\
        );

    \I__4032\ : InMux
    port map (
            O => \N__16842\,
            I => \N__16802\
        );

    \I__4031\ : InMux
    port map (
            O => \N__16841\,
            I => \N__16802\
        );

    \I__4030\ : InMux
    port map (
            O => \N__16840\,
            I => \N__16802\
        );

    \I__4029\ : InMux
    port map (
            O => \N__16837\,
            I => \N__16802\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__16826\,
            I => \N__16799\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__16821\,
            I => \Lab_UT_di_Mones_1\
        );

    \I__4026\ : Odrv4
    port map (
            O => \N__16816\,
            I => \Lab_UT_di_Mones_1\
        );

    \I__4025\ : LocalMux
    port map (
            O => \N__16813\,
            I => \Lab_UT_di_Mones_1\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__16802\,
            I => \Lab_UT_di_Mones_1\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__16799\,
            I => \Lab_UT_di_Mones_1\
        );

    \I__4022\ : CascadeMux
    port map (
            O => \N__16788\,
            I => \N__16785\
        );

    \I__4021\ : InMux
    port map (
            O => \N__16785\,
            I => \N__16777\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__16784\,
            I => \N__16774\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__16783\,
            I => \N__16771\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__16782\,
            I => \N__16768\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__16781\,
            I => \N__16764\
        );

    \I__4016\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16761\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__16777\,
            I => \N__16758\
        );

    \I__4014\ : InMux
    port map (
            O => \N__16774\,
            I => \N__16755\
        );

    \I__4013\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16751\
        );

    \I__4012\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16744\
        );

    \I__4011\ : InMux
    port map (
            O => \N__16767\,
            I => \N__16744\
        );

    \I__4010\ : InMux
    port map (
            O => \N__16764\,
            I => \N__16744\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__16761\,
            I => \N__16738\
        );

    \I__4008\ : Span4Mux_v
    port map (
            O => \N__16758\,
            I => \N__16733\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__16755\,
            I => \N__16733\
        );

    \I__4006\ : InMux
    port map (
            O => \N__16754\,
            I => \N__16730\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__16751\,
            I => \N__16725\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__16744\,
            I => \N__16725\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__16743\,
            I => \N__16722\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__16742\,
            I => \N__16717\
        );

    \I__4001\ : InMux
    port map (
            O => \N__16741\,
            I => \N__16713\
        );

    \I__4000\ : Span4Mux_v
    port map (
            O => \N__16738\,
            I => \N__16708\
        );

    \I__3999\ : Span4Mux_v
    port map (
            O => \N__16733\,
            I => \N__16708\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__16730\,
            I => \N__16703\
        );

    \I__3997\ : Span4Mux_h
    port map (
            O => \N__16725\,
            I => \N__16703\
        );

    \I__3996\ : InMux
    port map (
            O => \N__16722\,
            I => \N__16692\
        );

    \I__3995\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16692\
        );

    \I__3994\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16692\
        );

    \I__3993\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16692\
        );

    \I__3992\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16692\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__16713\,
            I => \Lab_UT_di_Mones_3\
        );

    \I__3990\ : Odrv4
    port map (
            O => \N__16708\,
            I => \Lab_UT_di_Mones_3\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__16703\,
            I => \Lab_UT_di_Mones_3\
        );

    \I__3988\ : LocalMux
    port map (
            O => \N__16692\,
            I => \Lab_UT_di_Mones_3\
        );

    \I__3987\ : InMux
    port map (
            O => \N__16683\,
            I => \N__16678\
        );

    \I__3986\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16675\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__16681\,
            I => \N__16665\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__16678\,
            I => \N__16662\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__16675\,
            I => \N__16653\
        );

    \I__3982\ : InMux
    port map (
            O => \N__16674\,
            I => \N__16642\
        );

    \I__3981\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16642\
        );

    \I__3980\ : InMux
    port map (
            O => \N__16672\,
            I => \N__16642\
        );

    \I__3979\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16642\
        );

    \I__3978\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16642\
        );

    \I__3977\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16639\
        );

    \I__3976\ : InMux
    port map (
            O => \N__16668\,
            I => \N__16636\
        );

    \I__3975\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16633\
        );

    \I__3974\ : Span4Mux_h
    port map (
            O => \N__16662\,
            I => \N__16630\
        );

    \I__3973\ : InMux
    port map (
            O => \N__16661\,
            I => \N__16627\
        );

    \I__3972\ : InMux
    port map (
            O => \N__16660\,
            I => \N__16616\
        );

    \I__3971\ : InMux
    port map (
            O => \N__16659\,
            I => \N__16616\
        );

    \I__3970\ : InMux
    port map (
            O => \N__16658\,
            I => \N__16616\
        );

    \I__3969\ : InMux
    port map (
            O => \N__16657\,
            I => \N__16616\
        );

    \I__3968\ : InMux
    port map (
            O => \N__16656\,
            I => \N__16616\
        );

    \I__3967\ : Span4Mux_h
    port map (
            O => \N__16653\,
            I => \N__16611\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__16642\,
            I => \N__16611\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__16639\,
            I => \Lab_UT_di_Mones_0\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__16636\,
            I => \Lab_UT_di_Mones_0\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__16633\,
            I => \Lab_UT_di_Mones_0\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__16630\,
            I => \Lab_UT_di_Mones_0\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__16627\,
            I => \Lab_UT_di_Mones_0\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__16616\,
            I => \Lab_UT_di_Mones_0\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__16611\,
            I => \Lab_UT_di_Mones_0\
        );

    \I__3958\ : InMux
    port map (
            O => \N__16596\,
            I => \N__16590\
        );

    \I__3957\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16590\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__16590\,
            I => \N__16587\
        );

    \I__3955\ : Span12Mux_s3_h
    port map (
            O => \N__16587\,
            I => \N__16584\
        );

    \I__3954\ : Odrv12
    port map (
            O => \N__16584\,
            I => \uu2.N_2160_1_0_0\
        );

    \I__3953\ : InMux
    port map (
            O => \N__16581\,
            I => \N__16578\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__16578\,
            I => \N__16574\
        );

    \I__3951\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16571\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__16574\,
            I => \N__16564\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__16571\,
            I => \N__16564\
        );

    \I__3948\ : InMux
    port map (
            O => \N__16570\,
            I => \N__16561\
        );

    \I__3947\ : InMux
    port map (
            O => \N__16569\,
            I => \N__16558\
        );

    \I__3946\ : Span4Mux_h
    port map (
            O => \N__16564\,
            I => \N__16553\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__16561\,
            I => \N__16553\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__16558\,
            I => \Lab_UT_dicRun\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__16553\,
            I => \Lab_UT_dicRun\
        );

    \I__3942\ : InMux
    port map (
            O => \N__16548\,
            I => \N__16543\
        );

    \I__3941\ : InMux
    port map (
            O => \N__16547\,
            I => \N__16538\
        );

    \I__3940\ : InMux
    port map (
            O => \N__16546\,
            I => \N__16534\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__16543\,
            I => \N__16531\
        );

    \I__3938\ : InMux
    port map (
            O => \N__16542\,
            I => \N__16526\
        );

    \I__3937\ : InMux
    port map (
            O => \N__16541\,
            I => \N__16526\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__16538\,
            I => \N__16523\
        );

    \I__3935\ : InMux
    port map (
            O => \N__16537\,
            I => \N__16520\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__16534\,
            I => \N__16517\
        );

    \I__3933\ : Span4Mux_v
    port map (
            O => \N__16531\,
            I => \N__16512\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__16526\,
            I => \N__16512\
        );

    \I__3931\ : Span4Mux_v
    port map (
            O => \N__16523\,
            I => \N__16509\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__16520\,
            I => \Lab_UT_l_oneSecPluse\
        );

    \I__3929\ : Odrv12
    port map (
            O => \N__16517\,
            I => \Lab_UT_l_oneSecPluse\
        );

    \I__3928\ : Odrv4
    port map (
            O => \N__16512\,
            I => \Lab_UT_l_oneSecPluse\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__16509\,
            I => \Lab_UT_l_oneSecPluse\
        );

    \I__3926\ : IoInMux
    port map (
            O => \N__16500\,
            I => \N__16497\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__16497\,
            I => \N__16494\
        );

    \I__3924\ : Odrv4
    port map (
            O => \N__16494\,
            I => led_c_4
        );

    \I__3923\ : InMux
    port map (
            O => \N__16491\,
            I => \N__16488\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__16488\,
            I => \uu2.un1_w_addr_displaying_46_1\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__16485\,
            I => \uu2.un1_w_addr_displaying_46_1_cascade_\
        );

    \I__3920\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16479\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__16479\,
            I => \N__16476\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__16476\,
            I => \uu2.w_addr_displaying_RNI8U3D2Z0Z_0\
        );

    \I__3917\ : InMux
    port map (
            O => \N__16473\,
            I => \N__16469\
        );

    \I__3916\ : InMux
    port map (
            O => \N__16472\,
            I => \N__16466\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__16469\,
            I => \N__16460\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__16466\,
            I => \N__16455\
        );

    \I__3913\ : InMux
    port map (
            O => \N__16465\,
            I => \N__16450\
        );

    \I__3912\ : InMux
    port map (
            O => \N__16464\,
            I => \N__16450\
        );

    \I__3911\ : InMux
    port map (
            O => \N__16463\,
            I => \N__16447\
        );

    \I__3910\ : Span4Mux_h
    port map (
            O => \N__16460\,
            I => \N__16444\
        );

    \I__3909\ : InMux
    port map (
            O => \N__16459\,
            I => \N__16441\
        );

    \I__3908\ : InMux
    port map (
            O => \N__16458\,
            I => \N__16438\
        );

    \I__3907\ : Span4Mux_h
    port map (
            O => \N__16455\,
            I => \N__16433\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__16450\,
            I => \N__16433\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__16447\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__16444\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__16441\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__16438\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__3901\ : Odrv4
    port map (
            O => \N__16433\,
            I => \uu2.w_addr_displaying_5_repZ0Z1\
        );

    \I__3900\ : InMux
    port map (
            O => \N__16422\,
            I => \N__16418\
        );

    \I__3899\ : InMux
    port map (
            O => \N__16421\,
            I => \N__16410\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__16418\,
            I => \N__16406\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__16417\,
            I => \N__16403\
        );

    \I__3896\ : InMux
    port map (
            O => \N__16416\,
            I => \N__16398\
        );

    \I__3895\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16398\
        );

    \I__3894\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16393\
        );

    \I__3893\ : InMux
    port map (
            O => \N__16413\,
            I => \N__16393\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__16410\,
            I => \N__16390\
        );

    \I__3891\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16387\
        );

    \I__3890\ : Span4Mux_h
    port map (
            O => \N__16406\,
            I => \N__16384\
        );

    \I__3889\ : InMux
    port map (
            O => \N__16403\,
            I => \N__16381\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__16398\,
            I => \N__16378\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__16393\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__3886\ : Odrv4
    port map (
            O => \N__16390\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__16387\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__16384\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__16381\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__16378\,
            I => \uu2.w_addr_displaying_6_repZ0Z1\
        );

    \I__3881\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16360\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__16364\,
            I => \N__16357\
        );

    \I__3879\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16354\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__16360\,
            I => \N__16351\
        );

    \I__3877\ : InMux
    port map (
            O => \N__16357\,
            I => \N__16348\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__16354\,
            I => \N__16337\
        );

    \I__3875\ : Span4Mux_h
    port map (
            O => \N__16351\,
            I => \N__16337\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__16348\,
            I => \N__16334\
        );

    \I__3873\ : InMux
    port map (
            O => \N__16347\,
            I => \N__16329\
        );

    \I__3872\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16329\
        );

    \I__3871\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16320\
        );

    \I__3870\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16320\
        );

    \I__3869\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16320\
        );

    \I__3868\ : InMux
    port map (
            O => \N__16342\,
            I => \N__16320\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__16337\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__3866\ : Odrv4
    port map (
            O => \N__16334\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__16329\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__16320\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__3863\ : InMux
    port map (
            O => \N__16311\,
            I => \N__16308\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__16308\,
            I => \uu2.un1_w_addr_displaying_38_1\
        );

    \I__3861\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16302\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__16302\,
            I => \N__16299\
        );

    \I__3859\ : Span4Mux_v
    port map (
            O => \N__16299\,
            I => \N__16296\
        );

    \I__3858\ : Odrv4
    port map (
            O => \N__16296\,
            I => \uu2.segment3_m_3Z0Z_1\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__16293\,
            I => \uu2.un1_w_addr_displaying_38_1_cascade_\
        );

    \I__3856\ : InMux
    port map (
            O => \N__16290\,
            I => \N__16280\
        );

    \I__3855\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16269\
        );

    \I__3854\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16269\
        );

    \I__3853\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16269\
        );

    \I__3852\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16269\
        );

    \I__3851\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16262\
        );

    \I__3850\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16262\
        );

    \I__3849\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16262\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__16280\,
            I => \N__16259\
        );

    \I__3847\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16254\
        );

    \I__3846\ : InMux
    port map (
            O => \N__16278\,
            I => \N__16254\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__16269\,
            I => \N__16248\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__16262\,
            I => \N__16245\
        );

    \I__3843\ : Span4Mux_h
    port map (
            O => \N__16259\,
            I => \N__16240\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__16254\,
            I => \N__16240\
        );

    \I__3841\ : InMux
    port map (
            O => \N__16253\,
            I => \N__16237\
        );

    \I__3840\ : InMux
    port map (
            O => \N__16252\,
            I => \N__16234\
        );

    \I__3839\ : InMux
    port map (
            O => \N__16251\,
            I => \N__16231\
        );

    \I__3838\ : Span4Mux_h
    port map (
            O => \N__16248\,
            I => \N__16228\
        );

    \I__3837\ : Span4Mux_v
    port map (
            O => \N__16245\,
            I => \N__16225\
        );

    \I__3836\ : Span4Mux_h
    port map (
            O => \N__16240\,
            I => \N__16218\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__16237\,
            I => \N__16218\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__16234\,
            I => \N__16218\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__16231\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__16228\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3831\ : Odrv4
    port map (
            O => \N__16225\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__16218\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3829\ : InMux
    port map (
            O => \N__16209\,
            I => \N__16206\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__16206\,
            I => \uu2.segment3_m_1\
        );

    \I__3827\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16194\
        );

    \I__3826\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16194\
        );

    \I__3825\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16188\
        );

    \I__3824\ : InMux
    port map (
            O => \N__16200\,
            I => \N__16188\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__16199\,
            I => \N__16185\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__16194\,
            I => \N__16180\
        );

    \I__3821\ : InMux
    port map (
            O => \N__16193\,
            I => \N__16177\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__16188\,
            I => \N__16172\
        );

    \I__3819\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16167\
        );

    \I__3818\ : InMux
    port map (
            O => \N__16184\,
            I => \N__16167\
        );

    \I__3817\ : InMux
    port map (
            O => \N__16183\,
            I => \N__16164\
        );

    \I__3816\ : Span4Mux_h
    port map (
            O => \N__16180\,
            I => \N__16161\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__16177\,
            I => \N__16158\
        );

    \I__3814\ : InMux
    port map (
            O => \N__16176\,
            I => \N__16153\
        );

    \I__3813\ : InMux
    port map (
            O => \N__16175\,
            I => \N__16153\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__16172\,
            I => \N__16147\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__16167\,
            I => \N__16147\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__16164\,
            I => \N__16144\
        );

    \I__3809\ : Span4Mux_v
    port map (
            O => \N__16161\,
            I => \N__16137\
        );

    \I__3808\ : Span4Mux_h
    port map (
            O => \N__16158\,
            I => \N__16137\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__16153\,
            I => \N__16137\
        );

    \I__3806\ : InMux
    port map (
            O => \N__16152\,
            I => \N__16131\
        );

    \I__3805\ : Span4Mux_h
    port map (
            O => \N__16147\,
            I => \N__16128\
        );

    \I__3804\ : Span12Mux_s11_v
    port map (
            O => \N__16144\,
            I => \N__16125\
        );

    \I__3803\ : Span4Mux_h
    port map (
            O => \N__16137\,
            I => \N__16122\
        );

    \I__3802\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16115\
        );

    \I__3801\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16115\
        );

    \I__3800\ : InMux
    port map (
            O => \N__16134\,
            I => \N__16115\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__16131\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__16128\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3797\ : Odrv12
    port map (
            O => \N__16125\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__16122\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__16115\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__16104\,
            I => \N__16099\
        );

    \I__3793\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16087\
        );

    \I__3792\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16084\
        );

    \I__3791\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16079\
        );

    \I__3790\ : InMux
    port map (
            O => \N__16098\,
            I => \N__16076\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__16097\,
            I => \N__16073\
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__16096\,
            I => \N__16070\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__16095\,
            I => \N__16067\
        );

    \I__3786\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16060\
        );

    \I__3785\ : InMux
    port map (
            O => \N__16093\,
            I => \N__16060\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__16092\,
            I => \N__16050\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__16091\,
            I => \N__16046\
        );

    \I__3782\ : InMux
    port map (
            O => \N__16090\,
            I => \N__16042\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__16087\,
            I => \N__16037\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__16084\,
            I => \N__16037\
        );

    \I__3779\ : InMux
    port map (
            O => \N__16083\,
            I => \N__16032\
        );

    \I__3778\ : InMux
    port map (
            O => \N__16082\,
            I => \N__16032\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__16079\,
            I => \N__16029\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__16076\,
            I => \N__16026\
        );

    \I__3775\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16023\
        );

    \I__3774\ : InMux
    port map (
            O => \N__16070\,
            I => \N__16014\
        );

    \I__3773\ : InMux
    port map (
            O => \N__16067\,
            I => \N__16014\
        );

    \I__3772\ : InMux
    port map (
            O => \N__16066\,
            I => \N__16014\
        );

    \I__3771\ : InMux
    port map (
            O => \N__16065\,
            I => \N__16014\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__16060\,
            I => \N__16011\
        );

    \I__3769\ : InMux
    port map (
            O => \N__16059\,
            I => \N__16006\
        );

    \I__3768\ : InMux
    port map (
            O => \N__16058\,
            I => \N__16006\
        );

    \I__3767\ : InMux
    port map (
            O => \N__16057\,
            I => \N__16001\
        );

    \I__3766\ : InMux
    port map (
            O => \N__16056\,
            I => \N__16001\
        );

    \I__3765\ : InMux
    port map (
            O => \N__16055\,
            I => \N__15994\
        );

    \I__3764\ : InMux
    port map (
            O => \N__16054\,
            I => \N__15994\
        );

    \I__3763\ : InMux
    port map (
            O => \N__16053\,
            I => \N__15994\
        );

    \I__3762\ : InMux
    port map (
            O => \N__16050\,
            I => \N__15989\
        );

    \I__3761\ : InMux
    port map (
            O => \N__16049\,
            I => \N__15989\
        );

    \I__3760\ : InMux
    port map (
            O => \N__16046\,
            I => \N__15984\
        );

    \I__3759\ : InMux
    port map (
            O => \N__16045\,
            I => \N__15984\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__16042\,
            I => \N__15981\
        );

    \I__3757\ : Span4Mux_v
    port map (
            O => \N__16037\,
            I => \N__15978\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__16032\,
            I => \N__15971\
        );

    \I__3755\ : Span4Mux_v
    port map (
            O => \N__16029\,
            I => \N__15971\
        );

    \I__3754\ : Span4Mux_h
    port map (
            O => \N__16026\,
            I => \N__15971\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__16023\,
            I => \N__15964\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__16014\,
            I => \N__15964\
        );

    \I__3751\ : Span4Mux_v
    port map (
            O => \N__16011\,
            I => \N__15964\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__16006\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__16001\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__15994\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__15989\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__15984\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__15981\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3744\ : Odrv4
    port map (
            O => \N__15978\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__15971\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__15964\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3741\ : InMux
    port map (
            O => \N__15945\,
            I => \N__15940\
        );

    \I__3740\ : InMux
    port map (
            O => \N__15944\,
            I => \N__15937\
        );

    \I__3739\ : InMux
    port map (
            O => \N__15943\,
            I => \N__15934\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__15940\,
            I => \N__15931\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__15937\,
            I => \N__15928\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__15934\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__3735\ : Odrv4
    port map (
            O => \N__15931\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__15928\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__3733\ : InMux
    port map (
            O => \N__15921\,
            I => \N__15914\
        );

    \I__3732\ : InMux
    port map (
            O => \N__15920\,
            I => \N__15911\
        );

    \I__3731\ : InMux
    port map (
            O => \N__15919\,
            I => \N__15906\
        );

    \I__3730\ : InMux
    port map (
            O => \N__15918\,
            I => \N__15906\
        );

    \I__3729\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15903\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__15914\,
            I => \N__15869\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__15911\,
            I => \N__15866\
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__15906\,
            I => \N__15863\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__15903\,
            I => \N__15860\
        );

    \I__3724\ : SRMux
    port map (
            O => \N__15902\,
            I => \N__15753\
        );

    \I__3723\ : SRMux
    port map (
            O => \N__15901\,
            I => \N__15753\
        );

    \I__3722\ : SRMux
    port map (
            O => \N__15900\,
            I => \N__15753\
        );

    \I__3721\ : SRMux
    port map (
            O => \N__15899\,
            I => \N__15753\
        );

    \I__3720\ : SRMux
    port map (
            O => \N__15898\,
            I => \N__15753\
        );

    \I__3719\ : SRMux
    port map (
            O => \N__15897\,
            I => \N__15753\
        );

    \I__3718\ : SRMux
    port map (
            O => \N__15896\,
            I => \N__15753\
        );

    \I__3717\ : SRMux
    port map (
            O => \N__15895\,
            I => \N__15753\
        );

    \I__3716\ : SRMux
    port map (
            O => \N__15894\,
            I => \N__15753\
        );

    \I__3715\ : SRMux
    port map (
            O => \N__15893\,
            I => \N__15753\
        );

    \I__3714\ : SRMux
    port map (
            O => \N__15892\,
            I => \N__15753\
        );

    \I__3713\ : SRMux
    port map (
            O => \N__15891\,
            I => \N__15753\
        );

    \I__3712\ : SRMux
    port map (
            O => \N__15890\,
            I => \N__15753\
        );

    \I__3711\ : SRMux
    port map (
            O => \N__15889\,
            I => \N__15753\
        );

    \I__3710\ : SRMux
    port map (
            O => \N__15888\,
            I => \N__15753\
        );

    \I__3709\ : SRMux
    port map (
            O => \N__15887\,
            I => \N__15753\
        );

    \I__3708\ : SRMux
    port map (
            O => \N__15886\,
            I => \N__15753\
        );

    \I__3707\ : SRMux
    port map (
            O => \N__15885\,
            I => \N__15753\
        );

    \I__3706\ : SRMux
    port map (
            O => \N__15884\,
            I => \N__15753\
        );

    \I__3705\ : SRMux
    port map (
            O => \N__15883\,
            I => \N__15753\
        );

    \I__3704\ : SRMux
    port map (
            O => \N__15882\,
            I => \N__15753\
        );

    \I__3703\ : SRMux
    port map (
            O => \N__15881\,
            I => \N__15753\
        );

    \I__3702\ : SRMux
    port map (
            O => \N__15880\,
            I => \N__15753\
        );

    \I__3701\ : SRMux
    port map (
            O => \N__15879\,
            I => \N__15753\
        );

    \I__3700\ : SRMux
    port map (
            O => \N__15878\,
            I => \N__15753\
        );

    \I__3699\ : SRMux
    port map (
            O => \N__15877\,
            I => \N__15753\
        );

    \I__3698\ : SRMux
    port map (
            O => \N__15876\,
            I => \N__15753\
        );

    \I__3697\ : SRMux
    port map (
            O => \N__15875\,
            I => \N__15753\
        );

    \I__3696\ : SRMux
    port map (
            O => \N__15874\,
            I => \N__15753\
        );

    \I__3695\ : SRMux
    port map (
            O => \N__15873\,
            I => \N__15753\
        );

    \I__3694\ : SRMux
    port map (
            O => \N__15872\,
            I => \N__15753\
        );

    \I__3693\ : Glb2LocalMux
    port map (
            O => \N__15869\,
            I => \N__15753\
        );

    \I__3692\ : Glb2LocalMux
    port map (
            O => \N__15866\,
            I => \N__15753\
        );

    \I__3691\ : Glb2LocalMux
    port map (
            O => \N__15863\,
            I => \N__15753\
        );

    \I__3690\ : Glb2LocalMux
    port map (
            O => \N__15860\,
            I => \N__15753\
        );

    \I__3689\ : SRMux
    port map (
            O => \N__15859\,
            I => \N__15753\
        );

    \I__3688\ : SRMux
    port map (
            O => \N__15858\,
            I => \N__15753\
        );

    \I__3687\ : SRMux
    port map (
            O => \N__15857\,
            I => \N__15753\
        );

    \I__3686\ : SRMux
    port map (
            O => \N__15856\,
            I => \N__15753\
        );

    \I__3685\ : SRMux
    port map (
            O => \N__15855\,
            I => \N__15753\
        );

    \I__3684\ : SRMux
    port map (
            O => \N__15854\,
            I => \N__15753\
        );

    \I__3683\ : SRMux
    port map (
            O => \N__15853\,
            I => \N__15753\
        );

    \I__3682\ : SRMux
    port map (
            O => \N__15852\,
            I => \N__15753\
        );

    \I__3681\ : SRMux
    port map (
            O => \N__15851\,
            I => \N__15753\
        );

    \I__3680\ : SRMux
    port map (
            O => \N__15850\,
            I => \N__15753\
        );

    \I__3679\ : SRMux
    port map (
            O => \N__15849\,
            I => \N__15753\
        );

    \I__3678\ : SRMux
    port map (
            O => \N__15848\,
            I => \N__15753\
        );

    \I__3677\ : GlobalMux
    port map (
            O => \N__15753\,
            I => \N__15750\
        );

    \I__3676\ : gio2CtrlBuf
    port map (
            O => \N__15750\,
            I => rst_g
        );

    \I__3675\ : InMux
    port map (
            O => \N__15747\,
            I => \N__15744\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__15744\,
            I => \N__15741\
        );

    \I__3673\ : Span4Mux_h
    port map (
            O => \N__15741\,
            I => \N__15738\
        );

    \I__3672\ : Odrv4
    port map (
            O => \N__15738\,
            I => \uu2.mem0.N_2160_2\
        );

    \I__3671\ : InMux
    port map (
            O => \N__15735\,
            I => \N__15726\
        );

    \I__3670\ : InMux
    port map (
            O => \N__15734\,
            I => \N__15716\
        );

    \I__3669\ : InMux
    port map (
            O => \N__15733\,
            I => \N__15716\
        );

    \I__3668\ : InMux
    port map (
            O => \N__15732\,
            I => \N__15716\
        );

    \I__3667\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15716\
        );

    \I__3666\ : InMux
    port map (
            O => \N__15730\,
            I => \N__15708\
        );

    \I__3665\ : InMux
    port map (
            O => \N__15729\,
            I => \N__15708\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__15726\,
            I => \N__15705\
        );

    \I__3663\ : InMux
    port map (
            O => \N__15725\,
            I => \N__15702\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__15716\,
            I => \N__15699\
        );

    \I__3661\ : InMux
    port map (
            O => \N__15715\,
            I => \N__15692\
        );

    \I__3660\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15692\
        );

    \I__3659\ : InMux
    port map (
            O => \N__15713\,
            I => \N__15692\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__15708\,
            I => \N__15686\
        );

    \I__3657\ : Span4Mux_v
    port map (
            O => \N__15705\,
            I => \N__15681\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__15702\,
            I => \N__15681\
        );

    \I__3655\ : Span12Mux_s9_v
    port map (
            O => \N__15699\,
            I => \N__15678\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__15692\,
            I => \N__15675\
        );

    \I__3653\ : InMux
    port map (
            O => \N__15691\,
            I => \N__15668\
        );

    \I__3652\ : InMux
    port map (
            O => \N__15690\,
            I => \N__15668\
        );

    \I__3651\ : InMux
    port map (
            O => \N__15689\,
            I => \N__15668\
        );

    \I__3650\ : Span4Mux_h
    port map (
            O => \N__15686\,
            I => \N__15665\
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__15681\,
            I => \Lab_UT_di_Sones_0\
        );

    \I__3648\ : Odrv12
    port map (
            O => \N__15678\,
            I => \Lab_UT_di_Sones_0\
        );

    \I__3647\ : Odrv12
    port map (
            O => \N__15675\,
            I => \Lab_UT_di_Sones_0\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__15668\,
            I => \Lab_UT_di_Sones_0\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__15665\,
            I => \Lab_UT_di_Sones_0\
        );

    \I__3644\ : InMux
    port map (
            O => \N__15654\,
            I => \N__15650\
        );

    \I__3643\ : InMux
    port map (
            O => \N__15653\,
            I => \N__15647\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__15650\,
            I => \N__15643\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__15647\,
            I => \N__15632\
        );

    \I__3640\ : InMux
    port map (
            O => \N__15646\,
            I => \N__15629\
        );

    \I__3639\ : Span4Mux_h
    port map (
            O => \N__15643\,
            I => \N__15623\
        );

    \I__3638\ : InMux
    port map (
            O => \N__15642\,
            I => \N__15620\
        );

    \I__3637\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15611\
        );

    \I__3636\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15611\
        );

    \I__3635\ : InMux
    port map (
            O => \N__15639\,
            I => \N__15611\
        );

    \I__3634\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15611\
        );

    \I__3633\ : InMux
    port map (
            O => \N__15637\,
            I => \N__15603\
        );

    \I__3632\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15603\
        );

    \I__3631\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15603\
        );

    \I__3630\ : Span4Mux_v
    port map (
            O => \N__15632\,
            I => \N__15598\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__15629\,
            I => \N__15598\
        );

    \I__3628\ : InMux
    port map (
            O => \N__15628\,
            I => \N__15591\
        );

    \I__3627\ : InMux
    port map (
            O => \N__15627\,
            I => \N__15591\
        );

    \I__3626\ : InMux
    port map (
            O => \N__15626\,
            I => \N__15591\
        );

    \I__3625\ : Sp12to4
    port map (
            O => \N__15623\,
            I => \N__15584\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__15620\,
            I => \N__15584\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__15611\,
            I => \N__15584\
        );

    \I__3622\ : InMux
    port map (
            O => \N__15610\,
            I => \N__15581\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__15603\,
            I => \Lab_UT_di_Stens_0\
        );

    \I__3620\ : Odrv4
    port map (
            O => \N__15598\,
            I => \Lab_UT_di_Stens_0\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__15591\,
            I => \Lab_UT_di_Stens_0\
        );

    \I__3618\ : Odrv12
    port map (
            O => \N__15584\,
            I => \Lab_UT_di_Stens_0\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__15581\,
            I => \Lab_UT_di_Stens_0\
        );

    \I__3616\ : InMux
    port map (
            O => \N__15570\,
            I => \N__15567\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__15567\,
            I => \uu2.w_addr_displaying_4_rep2_RNI4S6JZ0\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__15564\,
            I => \uu2.w_addr_displaying_fast_RNIEDBMZ0Z_7_cascade_\
        );

    \I__3613\ : InMux
    port map (
            O => \N__15561\,
            I => \N__15558\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__15558\,
            I => \N__15555\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__15555\,
            I => \uu2.un1_segment4_sn_N_38_0\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__15552\,
            I => \N__15548\
        );

    \I__3609\ : InMux
    port map (
            O => \N__15551\,
            I => \N__15540\
        );

    \I__3608\ : InMux
    port map (
            O => \N__15548\,
            I => \N__15540\
        );

    \I__3607\ : InMux
    port map (
            O => \N__15547\,
            I => \N__15537\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__15546\,
            I => \N__15534\
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__15545\,
            I => \N__15527\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__15540\,
            I => \N__15523\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__15537\,
            I => \N__15520\
        );

    \I__3602\ : InMux
    port map (
            O => \N__15534\,
            I => \N__15515\
        );

    \I__3601\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15515\
        );

    \I__3600\ : InMux
    port map (
            O => \N__15532\,
            I => \N__15510\
        );

    \I__3599\ : InMux
    port map (
            O => \N__15531\,
            I => \N__15510\
        );

    \I__3598\ : InMux
    port map (
            O => \N__15530\,
            I => \N__15503\
        );

    \I__3597\ : InMux
    port map (
            O => \N__15527\,
            I => \N__15503\
        );

    \I__3596\ : InMux
    port map (
            O => \N__15526\,
            I => \N__15503\
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__15523\,
            I => \uu2.w_addr_displaying_4_repZ0Z2\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__15520\,
            I => \uu2.w_addr_displaying_4_repZ0Z2\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__15515\,
            I => \uu2.w_addr_displaying_4_repZ0Z2\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__15510\,
            I => \uu2.w_addr_displaying_4_repZ0Z2\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__15503\,
            I => \uu2.w_addr_displaying_4_repZ0Z2\
        );

    \I__3590\ : InMux
    port map (
            O => \N__15492\,
            I => \N__15487\
        );

    \I__3589\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15484\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__15490\,
            I => \N__15481\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__15487\,
            I => \N__15477\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__15484\,
            I => \N__15474\
        );

    \I__3585\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15471\
        );

    \I__3584\ : InMux
    port map (
            O => \N__15480\,
            I => \N__15468\
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__15477\,
            I => \uu2.N_111\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__15474\,
            I => \uu2.N_111\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__15471\,
            I => \uu2.N_111\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__15468\,
            I => \uu2.N_111\
        );

    \I__3579\ : InMux
    port map (
            O => \N__15459\,
            I => \N__15453\
        );

    \I__3578\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15446\
        );

    \I__3577\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15443\
        );

    \I__3576\ : CascadeMux
    port map (
            O => \N__15456\,
            I => \N__15438\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__15453\,
            I => \N__15435\
        );

    \I__3574\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15432\
        );

    \I__3573\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15427\
        );

    \I__3572\ : InMux
    port map (
            O => \N__15450\,
            I => \N__15427\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__15449\,
            I => \N__15422\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__15446\,
            I => \N__15415\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__15443\,
            I => \N__15415\
        );

    \I__3568\ : InMux
    port map (
            O => \N__15442\,
            I => \N__15412\
        );

    \I__3567\ : InMux
    port map (
            O => \N__15441\,
            I => \N__15409\
        );

    \I__3566\ : InMux
    port map (
            O => \N__15438\,
            I => \N__15406\
        );

    \I__3565\ : Span4Mux_h
    port map (
            O => \N__15435\,
            I => \N__15403\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__15432\,
            I => \N__15398\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__15427\,
            I => \N__15398\
        );

    \I__3562\ : InMux
    port map (
            O => \N__15426\,
            I => \N__15393\
        );

    \I__3561\ : InMux
    port map (
            O => \N__15425\,
            I => \N__15393\
        );

    \I__3560\ : InMux
    port map (
            O => \N__15422\,
            I => \N__15386\
        );

    \I__3559\ : InMux
    port map (
            O => \N__15421\,
            I => \N__15386\
        );

    \I__3558\ : InMux
    port map (
            O => \N__15420\,
            I => \N__15386\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__15415\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__15412\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__15409\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__15406\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__15403\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__15398\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__15393\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__15386\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3549\ : InMux
    port map (
            O => \N__15369\,
            I => \N__15362\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__15368\,
            I => \N__15359\
        );

    \I__3547\ : InMux
    port map (
            O => \N__15367\,
            I => \N__15356\
        );

    \I__3546\ : InMux
    port map (
            O => \N__15366\,
            I => \N__15353\
        );

    \I__3545\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15350\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__15362\,
            I => \N__15347\
        );

    \I__3543\ : InMux
    port map (
            O => \N__15359\,
            I => \N__15342\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__15356\,
            I => \N__15339\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__15353\,
            I => \N__15334\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__15350\,
            I => \N__15334\
        );

    \I__3539\ : Span4Mux_v
    port map (
            O => \N__15347\,
            I => \N__15331\
        );

    \I__3538\ : InMux
    port map (
            O => \N__15346\,
            I => \N__15326\
        );

    \I__3537\ : InMux
    port map (
            O => \N__15345\,
            I => \N__15326\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__15342\,
            I => \N__15321\
        );

    \I__3535\ : Span4Mux_h
    port map (
            O => \N__15339\,
            I => \N__15321\
        );

    \I__3534\ : Span4Mux_v
    port map (
            O => \N__15334\,
            I => \N__15318\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__15331\,
            I => \uu2.Z_decfrac106_6\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__15326\,
            I => \uu2.Z_decfrac106_6\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__15321\,
            I => \uu2.Z_decfrac106_6\
        );

    \I__3530\ : Odrv4
    port map (
            O => \N__15318\,
            I => \uu2.Z_decfrac106_6\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__15309\,
            I => \N__15302\
        );

    \I__3528\ : InMux
    port map (
            O => \N__15308\,
            I => \N__15296\
        );

    \I__3527\ : InMux
    port map (
            O => \N__15307\,
            I => \N__15296\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__15306\,
            I => \N__15293\
        );

    \I__3525\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15288\
        );

    \I__3524\ : InMux
    port map (
            O => \N__15302\,
            I => \N__15283\
        );

    \I__3523\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15283\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__15296\,
            I => \N__15280\
        );

    \I__3521\ : InMux
    port map (
            O => \N__15293\,
            I => \N__15275\
        );

    \I__3520\ : InMux
    port map (
            O => \N__15292\,
            I => \N__15275\
        );

    \I__3519\ : InMux
    port map (
            O => \N__15291\,
            I => \N__15272\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__15288\,
            I => \N__15267\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__15283\,
            I => \N__15267\
        );

    \I__3516\ : Span4Mux_h
    port map (
            O => \N__15280\,
            I => \N__15264\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__15275\,
            I => \N__15261\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__15272\,
            I => \N__15256\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__15267\,
            I => \N__15256\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__15264\,
            I => \uu2.un15_w_data_displaying_5\
        );

    \I__3511\ : Odrv4
    port map (
            O => \N__15261\,
            I => \uu2.un15_w_data_displaying_5\
        );

    \I__3510\ : Odrv4
    port map (
            O => \N__15256\,
            I => \uu2.un15_w_data_displaying_5\
        );

    \I__3509\ : InMux
    port map (
            O => \N__15249\,
            I => \N__15244\
        );

    \I__3508\ : InMux
    port map (
            O => \N__15248\,
            I => \N__15241\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__15247\,
            I => \N__15237\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__15244\,
            I => \N__15232\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__15241\,
            I => \N__15229\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__15240\,
            I => \N__15226\
        );

    \I__3503\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15223\
        );

    \I__3502\ : InMux
    port map (
            O => \N__15236\,
            I => \N__15218\
        );

    \I__3501\ : InMux
    port map (
            O => \N__15235\,
            I => \N__15218\
        );

    \I__3500\ : Span4Mux_h
    port map (
            O => \N__15232\,
            I => \N__15215\
        );

    \I__3499\ : Span4Mux_h
    port map (
            O => \N__15229\,
            I => \N__15212\
        );

    \I__3498\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15209\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__15223\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__15218\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__15215\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__15212\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__15209\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__15198\,
            I => \L3_segment4_2_cascade_\
        );

    \I__3491\ : InMux
    port map (
            O => \N__15195\,
            I => \N__15192\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__15192\,
            I => \uu2.N_280\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__15189\,
            I => \N__15184\
        );

    \I__3488\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15179\
        );

    \I__3487\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15176\
        );

    \I__3486\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15173\
        );

    \I__3485\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15168\
        );

    \I__3484\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15168\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__15179\,
            I => \N__15163\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__15176\,
            I => \N__15160\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__15173\,
            I => \N__15157\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__15168\,
            I => \N__15154\
        );

    \I__3479\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15149\
        );

    \I__3478\ : InMux
    port map (
            O => \N__15166\,
            I => \N__15149\
        );

    \I__3477\ : Span4Mux_v
    port map (
            O => \N__15163\,
            I => \N__15138\
        );

    \I__3476\ : Span4Mux_h
    port map (
            O => \N__15160\,
            I => \N__15138\
        );

    \I__3475\ : Span4Mux_h
    port map (
            O => \N__15157\,
            I => \N__15138\
        );

    \I__3474\ : Span4Mux_h
    port map (
            O => \N__15154\,
            I => \N__15138\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__15149\,
            I => \N__15138\
        );

    \I__3472\ : Span4Mux_v
    port map (
            O => \N__15138\,
            I => \N__15127\
        );

    \I__3471\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15120\
        );

    \I__3470\ : InMux
    port map (
            O => \N__15136\,
            I => \N__15120\
        );

    \I__3469\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15120\
        );

    \I__3468\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15109\
        );

    \I__3467\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15109\
        );

    \I__3466\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15109\
        );

    \I__3465\ : InMux
    port map (
            O => \N__15131\,
            I => \N__15109\
        );

    \I__3464\ : InMux
    port map (
            O => \N__15130\,
            I => \N__15109\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__15127\,
            I => \Lab_UT_di_Mtens_2\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__15120\,
            I => \Lab_UT_di_Mtens_2\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__15109\,
            I => \Lab_UT_di_Mtens_2\
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__15102\,
            I => \N__15096\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__15101\,
            I => \N__15092\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__15100\,
            I => \N__15089\
        );

    \I__3457\ : InMux
    port map (
            O => \N__15099\,
            I => \N__15085\
        );

    \I__3456\ : InMux
    port map (
            O => \N__15096\,
            I => \N__15082\
        );

    \I__3455\ : InMux
    port map (
            O => \N__15095\,
            I => \N__15079\
        );

    \I__3454\ : InMux
    port map (
            O => \N__15092\,
            I => \N__15074\
        );

    \I__3453\ : InMux
    port map (
            O => \N__15089\,
            I => \N__15074\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__15088\,
            I => \N__15070\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__15085\,
            I => \N__15067\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__15082\,
            I => \N__15064\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__15079\,
            I => \N__15061\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__15074\,
            I => \N__15058\
        );

    \I__3447\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15053\
        );

    \I__3446\ : InMux
    port map (
            O => \N__15070\,
            I => \N__15053\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__15067\,
            I => \N__15043\
        );

    \I__3444\ : Span4Mux_h
    port map (
            O => \N__15064\,
            I => \N__15034\
        );

    \I__3443\ : Span4Mux_h
    port map (
            O => \N__15061\,
            I => \N__15034\
        );

    \I__3442\ : Span4Mux_h
    port map (
            O => \N__15058\,
            I => \N__15034\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__15053\,
            I => \N__15034\
        );

    \I__3440\ : InMux
    port map (
            O => \N__15052\,
            I => \N__15027\
        );

    \I__3439\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15027\
        );

    \I__3438\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15027\
        );

    \I__3437\ : InMux
    port map (
            O => \N__15049\,
            I => \N__15018\
        );

    \I__3436\ : InMux
    port map (
            O => \N__15048\,
            I => \N__15018\
        );

    \I__3435\ : InMux
    port map (
            O => \N__15047\,
            I => \N__15018\
        );

    \I__3434\ : InMux
    port map (
            O => \N__15046\,
            I => \N__15018\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__15043\,
            I => \Lab_UT_di_Mtens_3\
        );

    \I__3432\ : Odrv4
    port map (
            O => \N__15034\,
            I => \Lab_UT_di_Mtens_3\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__15027\,
            I => \Lab_UT_di_Mtens_3\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__15018\,
            I => \Lab_UT_di_Mtens_3\
        );

    \I__3429\ : InMux
    port map (
            O => \N__15009\,
            I => \N__15006\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__15006\,
            I => \L3_segment4_4\
        );

    \I__3427\ : InMux
    port map (
            O => \N__15003\,
            I => \N__14995\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__15002\,
            I => \N__14989\
        );

    \I__3425\ : InMux
    port map (
            O => \N__15001\,
            I => \N__14984\
        );

    \I__3424\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14979\
        );

    \I__3423\ : InMux
    port map (
            O => \N__14999\,
            I => \N__14979\
        );

    \I__3422\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14976\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__14995\,
            I => \N__14972\
        );

    \I__3420\ : InMux
    port map (
            O => \N__14994\,
            I => \N__14965\
        );

    \I__3419\ : InMux
    port map (
            O => \N__14993\,
            I => \N__14965\
        );

    \I__3418\ : InMux
    port map (
            O => \N__14992\,
            I => \N__14965\
        );

    \I__3417\ : InMux
    port map (
            O => \N__14989\,
            I => \N__14962\
        );

    \I__3416\ : InMux
    port map (
            O => \N__14988\,
            I => \N__14958\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__14987\,
            I => \N__14955\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__14984\,
            I => \N__14950\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__14979\,
            I => \N__14950\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__14976\,
            I => \N__14947\
        );

    \I__3411\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14944\
        );

    \I__3410\ : Span4Mux_v
    port map (
            O => \N__14972\,
            I => \N__14937\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__14965\,
            I => \N__14937\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__14962\,
            I => \N__14937\
        );

    \I__3407\ : InMux
    port map (
            O => \N__14961\,
            I => \N__14934\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__14958\,
            I => \N__14931\
        );

    \I__3405\ : InMux
    port map (
            O => \N__14955\,
            I => \N__14928\
        );

    \I__3404\ : Span4Mux_h
    port map (
            O => \N__14950\,
            I => \N__14925\
        );

    \I__3403\ : Span4Mux_h
    port map (
            O => \N__14947\,
            I => \N__14918\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__14944\,
            I => \N__14918\
        );

    \I__3401\ : Span4Mux_h
    port map (
            O => \N__14937\,
            I => \N__14918\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__14934\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__3399\ : Odrv4
    port map (
            O => \N__14931\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__14928\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__14925\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__14918\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__14907\,
            I => \N__14903\
        );

    \I__3394\ : InMux
    port map (
            O => \N__14906\,
            I => \N__14897\
        );

    \I__3393\ : InMux
    port map (
            O => \N__14903\,
            I => \N__14897\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__14902\,
            I => \N__14893\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__14897\,
            I => \N__14884\
        );

    \I__3390\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14881\
        );

    \I__3389\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14878\
        );

    \I__3388\ : InMux
    port map (
            O => \N__14892\,
            I => \N__14875\
        );

    \I__3387\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14870\
        );

    \I__3386\ : InMux
    port map (
            O => \N__14890\,
            I => \N__14870\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__14889\,
            I => \N__14867\
        );

    \I__3384\ : InMux
    port map (
            O => \N__14888\,
            I => \N__14861\
        );

    \I__3383\ : InMux
    port map (
            O => \N__14887\,
            I => \N__14861\
        );

    \I__3382\ : Span4Mux_v
    port map (
            O => \N__14884\,
            I => \N__14856\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__14881\,
            I => \N__14856\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__14878\,
            I => \N__14851\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__14875\,
            I => \N__14851\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__14870\,
            I => \N__14848\
        );

    \I__3377\ : InMux
    port map (
            O => \N__14867\,
            I => \N__14843\
        );

    \I__3376\ : InMux
    port map (
            O => \N__14866\,
            I => \N__14843\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__14861\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3374\ : Odrv4
    port map (
            O => \N__14856\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__14851\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__14848\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__14843\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3370\ : InMux
    port map (
            O => \N__14832\,
            I => \N__14828\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__14831\,
            I => \N__14823\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__14828\,
            I => \N__14817\
        );

    \I__3367\ : InMux
    port map (
            O => \N__14827\,
            I => \N__14814\
        );

    \I__3366\ : InMux
    port map (
            O => \N__14826\,
            I => \N__14809\
        );

    \I__3365\ : InMux
    port map (
            O => \N__14823\,
            I => \N__14809\
        );

    \I__3364\ : InMux
    port map (
            O => \N__14822\,
            I => \N__14806\
        );

    \I__3363\ : InMux
    port map (
            O => \N__14821\,
            I => \N__14801\
        );

    \I__3362\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14801\
        );

    \I__3361\ : Span4Mux_h
    port map (
            O => \N__14817\,
            I => \N__14796\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__14814\,
            I => \N__14796\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__14809\,
            I => \N__14793\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__14806\,
            I => \N__14787\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__14801\,
            I => \N__14780\
        );

    \I__3356\ : Span4Mux_h
    port map (
            O => \N__14796\,
            I => \N__14780\
        );

    \I__3355\ : Span4Mux_v
    port map (
            O => \N__14793\,
            I => \N__14780\
        );

    \I__3354\ : InMux
    port map (
            O => \N__14792\,
            I => \N__14773\
        );

    \I__3353\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14773\
        );

    \I__3352\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14773\
        );

    \I__3351\ : Odrv4
    port map (
            O => \N__14787\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__3350\ : Odrv4
    port map (
            O => \N__14780\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__14773\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__14766\,
            I => \N__14763\
        );

    \I__3347\ : InMux
    port map (
            O => \N__14763\,
            I => \N__14760\
        );

    \I__3346\ : LocalMux
    port map (
            O => \N__14760\,
            I => \N__14757\
        );

    \I__3345\ : Span4Mux_h
    port map (
            O => \N__14757\,
            I => \N__14754\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__14754\,
            I => \uu2.un1_segment3_m4_s_2_1\
        );

    \I__3343\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14738\
        );

    \I__3342\ : InMux
    port map (
            O => \N__14750\,
            I => \N__14738\
        );

    \I__3341\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14735\
        );

    \I__3340\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14721\
        );

    \I__3339\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14721\
        );

    \I__3338\ : InMux
    port map (
            O => \N__14746\,
            I => \N__14721\
        );

    \I__3337\ : InMux
    port map (
            O => \N__14745\,
            I => \N__14721\
        );

    \I__3336\ : InMux
    port map (
            O => \N__14744\,
            I => \N__14721\
        );

    \I__3335\ : InMux
    port map (
            O => \N__14743\,
            I => \N__14721\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__14738\,
            I => \N__14716\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__14735\,
            I => \N__14713\
        );

    \I__3332\ : InMux
    port map (
            O => \N__14734\,
            I => \N__14710\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__14721\,
            I => \N__14707\
        );

    \I__3330\ : InMux
    port map (
            O => \N__14720\,
            I => \N__14702\
        );

    \I__3329\ : InMux
    port map (
            O => \N__14719\,
            I => \N__14702\
        );

    \I__3328\ : Span4Mux_v
    port map (
            O => \N__14716\,
            I => \N__14699\
        );

    \I__3327\ : Span4Mux_s3_h
    port map (
            O => \N__14713\,
            I => \N__14696\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__14710\,
            I => \N__14693\
        );

    \I__3325\ : Span4Mux_v
    port map (
            O => \N__14707\,
            I => \N__14686\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__14702\,
            I => \N__14686\
        );

    \I__3323\ : Span4Mux_h
    port map (
            O => \N__14699\,
            I => \N__14686\
        );

    \I__3322\ : Odrv4
    port map (
            O => \N__14696\,
            I => \Lab_UT_di_Sones_2\
        );

    \I__3321\ : Odrv12
    port map (
            O => \N__14693\,
            I => \Lab_UT_di_Sones_2\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__14686\,
            I => \Lab_UT_di_Sones_2\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__14679\,
            I => \N__14676\
        );

    \I__3318\ : InMux
    port map (
            O => \N__14676\,
            I => \N__14668\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__14675\,
            I => \N__14665\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__14674\,
            I => \N__14661\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__14673\,
            I => \N__14658\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__14672\,
            I => \N__14655\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__14671\,
            I => \N__14652\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__14668\,
            I => \N__14647\
        );

    \I__3311\ : InMux
    port map (
            O => \N__14665\,
            I => \N__14638\
        );

    \I__3310\ : InMux
    port map (
            O => \N__14664\,
            I => \N__14638\
        );

    \I__3309\ : InMux
    port map (
            O => \N__14661\,
            I => \N__14638\
        );

    \I__3308\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14638\
        );

    \I__3307\ : InMux
    port map (
            O => \N__14655\,
            I => \N__14634\
        );

    \I__3306\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14629\
        );

    \I__3305\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14629\
        );

    \I__3304\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14626\
        );

    \I__3303\ : Span4Mux_h
    port map (
            O => \N__14647\,
            I => \N__14623\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__14638\,
            I => \N__14620\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__14637\,
            I => \N__14616\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__14634\,
            I => \N__14613\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__14629\,
            I => \N__14610\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__14626\,
            I => \N__14605\
        );

    \I__3297\ : Span4Mux_h
    port map (
            O => \N__14623\,
            I => \N__14605\
        );

    \I__3296\ : Span4Mux_h
    port map (
            O => \N__14620\,
            I => \N__14602\
        );

    \I__3295\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14597\
        );

    \I__3294\ : InMux
    port map (
            O => \N__14616\,
            I => \N__14597\
        );

    \I__3293\ : Span4Mux_v
    port map (
            O => \N__14613\,
            I => \N__14592\
        );

    \I__3292\ : Span4Mux_h
    port map (
            O => \N__14610\,
            I => \N__14592\
        );

    \I__3291\ : Sp12to4
    port map (
            O => \N__14605\,
            I => \N__14587\
        );

    \I__3290\ : Sp12to4
    port map (
            O => \N__14602\,
            I => \N__14587\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__14597\,
            I => \Lab_UT_di_Sones_3\
        );

    \I__3288\ : Odrv4
    port map (
            O => \N__14592\,
            I => \Lab_UT_di_Sones_3\
        );

    \I__3287\ : Odrv12
    port map (
            O => \N__14587\,
            I => \Lab_UT_di_Sones_3\
        );

    \I__3286\ : InMux
    port map (
            O => \N__14580\,
            I => \N__14577\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__14577\,
            I => \uu2.un1_segment3_m0\
        );

    \I__3284\ : InMux
    port map (
            O => \N__14574\,
            I => \N__14569\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__14573\,
            I => \N__14565\
        );

    \I__3282\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14562\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__14569\,
            I => \N__14559\
        );

    \I__3280\ : InMux
    port map (
            O => \N__14568\,
            I => \N__14551\
        );

    \I__3279\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14548\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__14562\,
            I => \N__14545\
        );

    \I__3277\ : Span4Mux_v
    port map (
            O => \N__14559\,
            I => \N__14542\
        );

    \I__3276\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14537\
        );

    \I__3275\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14537\
        );

    \I__3274\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14530\
        );

    \I__3273\ : InMux
    port map (
            O => \N__14555\,
            I => \N__14530\
        );

    \I__3272\ : InMux
    port map (
            O => \N__14554\,
            I => \N__14530\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__14551\,
            I => \N__14527\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__14548\,
            I => \uu2.w_addr_displaying_fastZ0Z_6\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__14545\,
            I => \uu2.w_addr_displaying_fastZ0Z_6\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__14542\,
            I => \uu2.w_addr_displaying_fastZ0Z_6\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__14537\,
            I => \uu2.w_addr_displaying_fastZ0Z_6\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__14530\,
            I => \uu2.w_addr_displaying_fastZ0Z_6\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__14527\,
            I => \uu2.w_addr_displaying_fastZ0Z_6\
        );

    \I__3264\ : CascadeMux
    port map (
            O => \N__14514\,
            I => \L3_segment1_3_cascade_\
        );

    \I__3263\ : InMux
    port map (
            O => \N__14511\,
            I => \N__14507\
        );

    \I__3262\ : InMux
    port map (
            O => \N__14510\,
            I => \N__14504\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__14507\,
            I => \N__14497\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__14504\,
            I => \N__14494\
        );

    \I__3259\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14491\
        );

    \I__3258\ : InMux
    port map (
            O => \N__14502\,
            I => \N__14484\
        );

    \I__3257\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14484\
        );

    \I__3256\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14484\
        );

    \I__3255\ : Span4Mux_h
    port map (
            O => \N__14497\,
            I => \N__14481\
        );

    \I__3254\ : Odrv4
    port map (
            O => \N__14494\,
            I => \uu2.w_addr_displaying_fastZ0Z_5\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__14491\,
            I => \uu2.w_addr_displaying_fastZ0Z_5\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__14484\,
            I => \uu2.w_addr_displaying_fastZ0Z_5\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__14481\,
            I => \uu2.w_addr_displaying_fastZ0Z_5\
        );

    \I__3250\ : InMux
    port map (
            O => \N__14472\,
            I => \N__14469\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__14469\,
            I => \N__14466\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__14466\,
            I => \uu2.w_addr_displaying_fast_RNIQD7R4Z0Z_5\
        );

    \I__3247\ : InMux
    port map (
            O => \N__14463\,
            I => \N__14458\
        );

    \I__3246\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14455\
        );

    \I__3245\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14450\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__14458\,
            I => \N__14447\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__14455\,
            I => \N__14444\
        );

    \I__3242\ : InMux
    port map (
            O => \N__14454\,
            I => \N__14439\
        );

    \I__3241\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14439\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__14450\,
            I => \N__14434\
        );

    \I__3239\ : Span4Mux_h
    port map (
            O => \N__14447\,
            I => \N__14434\
        );

    \I__3238\ : Odrv4
    port map (
            O => \N__14444\,
            I => \uu2.N_315_1\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__14439\,
            I => \uu2.N_315_1\
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__14434\,
            I => \uu2.N_315_1\
        );

    \I__3235\ : InMux
    port map (
            O => \N__14427\,
            I => \N__14422\
        );

    \I__3234\ : InMux
    port map (
            O => \N__14426\,
            I => \N__14417\
        );

    \I__3233\ : InMux
    port map (
            O => \N__14425\,
            I => \N__14417\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__14422\,
            I => \N__14410\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__14417\,
            I => \N__14410\
        );

    \I__3230\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14405\
        );

    \I__3229\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14405\
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__14410\,
            I => \uu2.w_addr_displaying_4_rep2_RNI75VMZ0\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__14405\,
            I => \uu2.w_addr_displaying_4_rep2_RNI75VMZ0\
        );

    \I__3226\ : InMux
    port map (
            O => \N__14400\,
            I => \N__14392\
        );

    \I__3225\ : InMux
    port map (
            O => \N__14399\,
            I => \N__14392\
        );

    \I__3224\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14387\
        );

    \I__3223\ : InMux
    port map (
            O => \N__14397\,
            I => \N__14387\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__14392\,
            I => \N__14381\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__14387\,
            I => \N__14378\
        );

    \I__3220\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14373\
        );

    \I__3219\ : InMux
    port map (
            O => \N__14385\,
            I => \N__14373\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__14384\,
            I => \N__14370\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__14381\,
            I => \N__14366\
        );

    \I__3216\ : Span4Mux_h
    port map (
            O => \N__14378\,
            I => \N__14363\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__14373\,
            I => \N__14360\
        );

    \I__3214\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14355\
        );

    \I__3213\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14355\
        );

    \I__3212\ : Odrv4
    port map (
            O => \N__14366\,
            I => \uu2.un1_segment3_m5\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__14363\,
            I => \uu2.un1_segment3_m5\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__14360\,
            I => \uu2.un1_segment3_m5\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__14355\,
            I => \uu2.un1_segment3_m5\
        );

    \I__3208\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14343\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__14343\,
            I => \uu2.N_813_0\
        );

    \I__3206\ : InMux
    port map (
            O => \N__14340\,
            I => \N__14337\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__14337\,
            I => \N__14334\
        );

    \I__3204\ : Odrv12
    port map (
            O => \N__14334\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_59\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__14331\,
            I => \N__14328\
        );

    \I__3202\ : InMux
    port map (
            O => \N__14328\,
            I => \N__14325\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__14325\,
            I => \N__14322\
        );

    \I__3200\ : Odrv12
    port map (
            O => \N__14322\,
            I => \uu2.segment2_m_2Z0Z_5\
        );

    \I__3199\ : InMux
    port map (
            O => \N__14319\,
            I => \N__14316\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__14316\,
            I => \uu2.segment2_m_5\
        );

    \I__3197\ : InMux
    port map (
            O => \N__14313\,
            I => \N__14309\
        );

    \I__3196\ : InMux
    port map (
            O => \N__14312\,
            I => \N__14303\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__14309\,
            I => \N__14300\
        );

    \I__3194\ : InMux
    port map (
            O => \N__14308\,
            I => \N__14295\
        );

    \I__3193\ : InMux
    port map (
            O => \N__14307\,
            I => \N__14295\
        );

    \I__3192\ : InMux
    port map (
            O => \N__14306\,
            I => \N__14292\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__14303\,
            I => \N__14289\
        );

    \I__3190\ : Span4Mux_h
    port map (
            O => \N__14300\,
            I => \N__14279\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__14295\,
            I => \N__14279\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__14292\,
            I => \N__14274\
        );

    \I__3187\ : Span4Mux_h
    port map (
            O => \N__14289\,
            I => \N__14274\
        );

    \I__3186\ : InMux
    port map (
            O => \N__14288\,
            I => \N__14271\
        );

    \I__3185\ : InMux
    port map (
            O => \N__14287\,
            I => \N__14262\
        );

    \I__3184\ : InMux
    port map (
            O => \N__14286\,
            I => \N__14262\
        );

    \I__3183\ : InMux
    port map (
            O => \N__14285\,
            I => \N__14262\
        );

    \I__3182\ : InMux
    port map (
            O => \N__14284\,
            I => \N__14262\
        );

    \I__3181\ : Odrv4
    port map (
            O => \N__14279\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3180\ : Odrv4
    port map (
            O => \N__14274\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__14271\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__14262\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3177\ : InMux
    port map (
            O => \N__14253\,
            I => \N__14250\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__14250\,
            I => \N__14247\
        );

    \I__3175\ : Span4Mux_v
    port map (
            O => \N__14247\,
            I => \N__14243\
        );

    \I__3174\ : InMux
    port map (
            O => \N__14246\,
            I => \N__14240\
        );

    \I__3173\ : Span4Mux_h
    port map (
            O => \N__14243\,
            I => \N__14235\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__14240\,
            I => \N__14235\
        );

    \I__3171\ : Span4Mux_v
    port map (
            O => \N__14235\,
            I => \N__14230\
        );

    \I__3170\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14227\
        );

    \I__3169\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14224\
        );

    \I__3168\ : Span4Mux_h
    port map (
            O => \N__14230\,
            I => \N__14214\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__14227\,
            I => \N__14214\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__14224\,
            I => \N__14214\
        );

    \I__3165\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14209\
        );

    \I__3164\ : InMux
    port map (
            O => \N__14222\,
            I => \N__14209\
        );

    \I__3163\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14206\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__14214\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__14209\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__14206\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3159\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14195\
        );

    \I__3158\ : InMux
    port map (
            O => \N__14198\,
            I => \N__14192\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__14195\,
            I => \N__14184\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__14192\,
            I => \N__14181\
        );

    \I__3155\ : InMux
    port map (
            O => \N__14191\,
            I => \N__14178\
        );

    \I__3154\ : InMux
    port map (
            O => \N__14190\,
            I => \N__14171\
        );

    \I__3153\ : InMux
    port map (
            O => \N__14189\,
            I => \N__14171\
        );

    \I__3152\ : InMux
    port map (
            O => \N__14188\,
            I => \N__14171\
        );

    \I__3151\ : InMux
    port map (
            O => \N__14187\,
            I => \N__14168\
        );

    \I__3150\ : Span4Mux_v
    port map (
            O => \N__14184\,
            I => \N__14162\
        );

    \I__3149\ : Span4Mux_v
    port map (
            O => \N__14181\,
            I => \N__14162\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__14178\,
            I => \N__14155\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__14171\,
            I => \N__14150\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__14168\,
            I => \N__14150\
        );

    \I__3145\ : InMux
    port map (
            O => \N__14167\,
            I => \N__14147\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__14162\,
            I => \N__14144\
        );

    \I__3143\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14135\
        );

    \I__3142\ : InMux
    port map (
            O => \N__14160\,
            I => \N__14135\
        );

    \I__3141\ : InMux
    port map (
            O => \N__14159\,
            I => \N__14135\
        );

    \I__3140\ : InMux
    port map (
            O => \N__14158\,
            I => \N__14135\
        );

    \I__3139\ : Span4Mux_h
    port map (
            O => \N__14155\,
            I => \N__14130\
        );

    \I__3138\ : Span4Mux_v
    port map (
            O => \N__14150\,
            I => \N__14130\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__14147\,
            I => \Lab_UT_di_Stens_2\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__14144\,
            I => \Lab_UT_di_Stens_2\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__14135\,
            I => \Lab_UT_di_Stens_2\
        );

    \I__3134\ : Odrv4
    port map (
            O => \N__14130\,
            I => \Lab_UT_di_Stens_2\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__14121\,
            I => \N__14117\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__14120\,
            I => \N__14114\
        );

    \I__3131\ : InMux
    port map (
            O => \N__14117\,
            I => \N__14107\
        );

    \I__3130\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14104\
        );

    \I__3129\ : CascadeMux
    port map (
            O => \N__14113\,
            I => \N__14101\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__14112\,
            I => \N__14098\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__14111\,
            I => \N__14095\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__14110\,
            I => \N__14092\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__14107\,
            I => \N__14083\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__14104\,
            I => \N__14083\
        );

    \I__3123\ : InMux
    port map (
            O => \N__14101\,
            I => \N__14080\
        );

    \I__3122\ : InMux
    port map (
            O => \N__14098\,
            I => \N__14075\
        );

    \I__3121\ : InMux
    port map (
            O => \N__14095\,
            I => \N__14075\
        );

    \I__3120\ : InMux
    port map (
            O => \N__14092\,
            I => \N__14072\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__14091\,
            I => \N__14067\
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__14090\,
            I => \N__14064\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__14089\,
            I => \N__14061\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__14088\,
            I => \N__14058\
        );

    \I__3115\ : Span4Mux_v
    port map (
            O => \N__14083\,
            I => \N__14055\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__14080\,
            I => \N__14048\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__14075\,
            I => \N__14048\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__14072\,
            I => \N__14048\
        );

    \I__3111\ : InMux
    port map (
            O => \N__14071\,
            I => \N__14043\
        );

    \I__3110\ : InMux
    port map (
            O => \N__14070\,
            I => \N__14043\
        );

    \I__3109\ : InMux
    port map (
            O => \N__14067\,
            I => \N__14036\
        );

    \I__3108\ : InMux
    port map (
            O => \N__14064\,
            I => \N__14036\
        );

    \I__3107\ : InMux
    port map (
            O => \N__14061\,
            I => \N__14036\
        );

    \I__3106\ : InMux
    port map (
            O => \N__14058\,
            I => \N__14033\
        );

    \I__3105\ : Span4Mux_h
    port map (
            O => \N__14055\,
            I => \N__14028\
        );

    \I__3104\ : Span4Mux_v
    port map (
            O => \N__14048\,
            I => \N__14028\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__14043\,
            I => \Lab_UT_di_Stens_3\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__14036\,
            I => \Lab_UT_di_Stens_3\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__14033\,
            I => \Lab_UT_di_Stens_3\
        );

    \I__3100\ : Odrv4
    port map (
            O => \N__14028\,
            I => \Lab_UT_di_Stens_3\
        );

    \I__3099\ : InMux
    port map (
            O => \N__14019\,
            I => \N__14016\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__14016\,
            I => \uu2.un1_segment3_m5_amZ0\
        );

    \I__3097\ : InMux
    port map (
            O => \N__14013\,
            I => \N__14007\
        );

    \I__3096\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14004\
        );

    \I__3095\ : InMux
    port map (
            O => \N__14011\,
            I => \N__14001\
        );

    \I__3094\ : InMux
    port map (
            O => \N__14010\,
            I => \N__13998\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__14007\,
            I => \N__13990\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__14004\,
            I => \N__13990\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__14001\,
            I => \N__13987\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__13998\,
            I => \N__13984\
        );

    \I__3089\ : InMux
    port map (
            O => \N__13997\,
            I => \N__13980\
        );

    \I__3088\ : InMux
    port map (
            O => \N__13996\,
            I => \N__13977\
        );

    \I__3087\ : InMux
    port map (
            O => \N__13995\,
            I => \N__13974\
        );

    \I__3086\ : Span4Mux_v
    port map (
            O => \N__13990\,
            I => \N__13969\
        );

    \I__3085\ : Span4Mux_v
    port map (
            O => \N__13987\,
            I => \N__13966\
        );

    \I__3084\ : Span4Mux_h
    port map (
            O => \N__13984\,
            I => \N__13963\
        );

    \I__3083\ : InMux
    port map (
            O => \N__13983\,
            I => \N__13960\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__13980\,
            I => \N__13957\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__13977\,
            I => \N__13952\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__13974\,
            I => \N__13952\
        );

    \I__3079\ : InMux
    port map (
            O => \N__13973\,
            I => \N__13949\
        );

    \I__3078\ : InMux
    port map (
            O => \N__13972\,
            I => \N__13946\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__13969\,
            I => \uu2.N_290_0_i_0\
        );

    \I__3076\ : Odrv4
    port map (
            O => \N__13966\,
            I => \uu2.N_290_0_i_0\
        );

    \I__3075\ : Odrv4
    port map (
            O => \N__13963\,
            I => \uu2.N_290_0_i_0\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__13960\,
            I => \uu2.N_290_0_i_0\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__13957\,
            I => \uu2.N_290_0_i_0\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__13952\,
            I => \uu2.N_290_0_i_0\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__13949\,
            I => \uu2.N_290_0_i_0\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__13946\,
            I => \uu2.N_290_0_i_0\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__13929\,
            I => \N__13926\
        );

    \I__3068\ : InMux
    port map (
            O => \N__13926\,
            I => \N__13920\
        );

    \I__3067\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13920\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__13920\,
            I => \N__13910\
        );

    \I__3065\ : InMux
    port map (
            O => \N__13919\,
            I => \N__13903\
        );

    \I__3064\ : InMux
    port map (
            O => \N__13918\,
            I => \N__13903\
        );

    \I__3063\ : InMux
    port map (
            O => \N__13917\,
            I => \N__13903\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__13916\,
            I => \N__13900\
        );

    \I__3061\ : InMux
    port map (
            O => \N__13915\,
            I => \N__13895\
        );

    \I__3060\ : InMux
    port map (
            O => \N__13914\,
            I => \N__13895\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__13913\,
            I => \N__13892\
        );

    \I__3058\ : Span4Mux_h
    port map (
            O => \N__13910\,
            I => \N__13889\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__13903\,
            I => \N__13886\
        );

    \I__3056\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13883\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__13895\,
            I => \N__13880\
        );

    \I__3054\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13877\
        );

    \I__3053\ : Sp12to4
    port map (
            O => \N__13889\,
            I => \N__13874\
        );

    \I__3052\ : Span4Mux_v
    port map (
            O => \N__13886\,
            I => \N__13871\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__13883\,
            I => \N__13866\
        );

    \I__3050\ : Span4Mux_h
    port map (
            O => \N__13880\,
            I => \N__13866\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__13877\,
            I => \uu2.un436_ci\
        );

    \I__3048\ : Odrv12
    port map (
            O => \N__13874\,
            I => \uu2.un436_ci\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__13871\,
            I => \uu2.un436_ci\
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__13866\,
            I => \uu2.un436_ci\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__13857\,
            I => \N__13853\
        );

    \I__3044\ : InMux
    port map (
            O => \N__13856\,
            I => \N__13848\
        );

    \I__3043\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13844\
        );

    \I__3042\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13838\
        );

    \I__3041\ : InMux
    port map (
            O => \N__13851\,
            I => \N__13838\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__13848\,
            I => \N__13835\
        );

    \I__3039\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13832\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__13844\,
            I => \N__13829\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__13843\,
            I => \N__13823\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__13838\,
            I => \N__13813\
        );

    \I__3035\ : Span4Mux_v
    port map (
            O => \N__13835\,
            I => \N__13813\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__13832\,
            I => \N__13813\
        );

    \I__3033\ : Span4Mux_s3_h
    port map (
            O => \N__13829\,
            I => \N__13813\
        );

    \I__3032\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13808\
        );

    \I__3031\ : InMux
    port map (
            O => \N__13827\,
            I => \N__13808\
        );

    \I__3030\ : InMux
    port map (
            O => \N__13826\,
            I => \N__13805\
        );

    \I__3029\ : InMux
    port map (
            O => \N__13823\,
            I => \N__13800\
        );

    \I__3028\ : InMux
    port map (
            O => \N__13822\,
            I => \N__13800\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__13813\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__13808\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__13805\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__13800\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__3023\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13788\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__13788\,
            I => \N__13785\
        );

    \I__3021\ : Odrv12
    port map (
            O => \N__13785\,
            I => \uu2.un1_w_addr_displaying_35_0\
        );

    \I__3020\ : InMux
    port map (
            O => \N__13782\,
            I => \N__13776\
        );

    \I__3019\ : InMux
    port map (
            O => \N__13781\,
            I => \N__13772\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__13780\,
            I => \N__13766\
        );

    \I__3017\ : InMux
    port map (
            O => \N__13779\,
            I => \N__13759\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__13776\,
            I => \N__13753\
        );

    \I__3015\ : InMux
    port map (
            O => \N__13775\,
            I => \N__13750\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__13772\,
            I => \N__13747\
        );

    \I__3013\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13744\
        );

    \I__3012\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13737\
        );

    \I__3011\ : InMux
    port map (
            O => \N__13769\,
            I => \N__13737\
        );

    \I__3010\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13737\
        );

    \I__3009\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13732\
        );

    \I__3008\ : InMux
    port map (
            O => \N__13764\,
            I => \N__13732\
        );

    \I__3007\ : InMux
    port map (
            O => \N__13763\,
            I => \N__13729\
        );

    \I__3006\ : InMux
    port map (
            O => \N__13762\,
            I => \N__13726\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__13759\,
            I => \N__13723\
        );

    \I__3004\ : InMux
    port map (
            O => \N__13758\,
            I => \N__13718\
        );

    \I__3003\ : InMux
    port map (
            O => \N__13757\,
            I => \N__13718\
        );

    \I__3002\ : InMux
    port map (
            O => \N__13756\,
            I => \N__13715\
        );

    \I__3001\ : Span4Mux_h
    port map (
            O => \N__13753\,
            I => \N__13708\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__13750\,
            I => \N__13708\
        );

    \I__2999\ : Span4Mux_h
    port map (
            O => \N__13747\,
            I => \N__13708\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__13744\,
            I => \N__13705\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__13737\,
            I => \N__13694\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__13732\,
            I => \N__13694\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__13729\,
            I => \N__13694\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__13726\,
            I => \N__13694\
        );

    \I__2993\ : Span4Mux_h
    port map (
            O => \N__13723\,
            I => \N__13694\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__13718\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__13715\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__13708\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__13705\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__13694\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__13683\,
            I => \uu2.un1_w_addr_displaying_35_0_cascade_\
        );

    \I__2986\ : InMux
    port map (
            O => \N__13680\,
            I => \N__13676\
        );

    \I__2985\ : InMux
    port map (
            O => \N__13679\,
            I => \N__13673\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__13676\,
            I => \uu2.un1_w_addr_displaying_inv_2\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__13673\,
            I => \uu2.un1_w_addr_displaying_inv_2\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__13668\,
            I => \uu2.N_813_0_cascade_\
        );

    \I__2981\ : InMux
    port map (
            O => \N__13665\,
            I => \N__13662\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__13662\,
            I => \N__13659\
        );

    \I__2979\ : Odrv12
    port map (
            O => \N__13659\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_58\
        );

    \I__2978\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13649\
        );

    \I__2977\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13649\
        );

    \I__2976\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13646\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__13649\,
            I => \N__13641\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__13646\,
            I => \N__13641\
        );

    \I__2973\ : Odrv12
    port map (
            O => \N__13641\,
            I => \Lab_UT.didpuu0.countEnMones\
        );

    \I__2972\ : InMux
    port map (
            O => \N__13638\,
            I => \N__13635\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__13635\,
            I => \N__13632\
        );

    \I__2970\ : Span4Mux_v
    port map (
            O => \N__13632\,
            I => \N__13629\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__13629\,
            I => \uu2.un1_segment3_m5_bmZ0\
        );

    \I__2968\ : InMux
    port map (
            O => \N__13626\,
            I => \N__13623\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__13623\,
            I => \N__13619\
        );

    \I__2966\ : InMux
    port map (
            O => \N__13622\,
            I => \N__13616\
        );

    \I__2965\ : Span4Mux_v
    port map (
            O => \N__13619\,
            I => \N__13612\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__13616\,
            I => \N__13609\
        );

    \I__2963\ : InMux
    port map (
            O => \N__13615\,
            I => \N__13606\
        );

    \I__2962\ : Odrv4
    port map (
            O => \N__13612\,
            I => bu_rx_data_1
        );

    \I__2961\ : Odrv12
    port map (
            O => \N__13609\,
            I => bu_rx_data_1
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__13606\,
            I => bu_rx_data_1
        );

    \I__2959\ : InMux
    port map (
            O => \N__13599\,
            I => \N__13596\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__13596\,
            I => \N__13593\
        );

    \I__2957\ : Sp12to4
    port map (
            O => \N__13593\,
            I => \N__13589\
        );

    \I__2956\ : InMux
    port map (
            O => \N__13592\,
            I => \N__13586\
        );

    \I__2955\ : Span12Mux_s11_v
    port map (
            O => \N__13589\,
            I => \N__13581\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__13586\,
            I => \N__13581\
        );

    \I__2953\ : Odrv12
    port map (
            O => \N__13581\,
            I => bu_rx_data_0
        );

    \I__2952\ : CEMux
    port map (
            O => \N__13578\,
            I => \N__13574\
        );

    \I__2951\ : CEMux
    port map (
            O => \N__13577\,
            I => \N__13571\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__13574\,
            I => \N__13567\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__13571\,
            I => \N__13564\
        );

    \I__2948\ : CEMux
    port map (
            O => \N__13570\,
            I => \N__13561\
        );

    \I__2947\ : Span4Mux_h
    port map (
            O => \N__13567\,
            I => \N__13554\
        );

    \I__2946\ : Span4Mux_h
    port map (
            O => \N__13564\,
            I => \N__13554\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__13561\,
            I => \N__13554\
        );

    \I__2944\ : Span4Mux_h
    port map (
            O => \N__13554\,
            I => \N__13551\
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__13551\,
            I => \buart.Z_rx.N_41_i\
        );

    \I__2942\ : ClkMux
    port map (
            O => \N__13548\,
            I => \N__13350\
        );

    \I__2941\ : ClkMux
    port map (
            O => \N__13547\,
            I => \N__13350\
        );

    \I__2940\ : ClkMux
    port map (
            O => \N__13546\,
            I => \N__13350\
        );

    \I__2939\ : ClkMux
    port map (
            O => \N__13545\,
            I => \N__13350\
        );

    \I__2938\ : ClkMux
    port map (
            O => \N__13544\,
            I => \N__13350\
        );

    \I__2937\ : ClkMux
    port map (
            O => \N__13543\,
            I => \N__13350\
        );

    \I__2936\ : ClkMux
    port map (
            O => \N__13542\,
            I => \N__13350\
        );

    \I__2935\ : ClkMux
    port map (
            O => \N__13541\,
            I => \N__13350\
        );

    \I__2934\ : ClkMux
    port map (
            O => \N__13540\,
            I => \N__13350\
        );

    \I__2933\ : ClkMux
    port map (
            O => \N__13539\,
            I => \N__13350\
        );

    \I__2932\ : ClkMux
    port map (
            O => \N__13538\,
            I => \N__13350\
        );

    \I__2931\ : ClkMux
    port map (
            O => \N__13537\,
            I => \N__13350\
        );

    \I__2930\ : ClkMux
    port map (
            O => \N__13536\,
            I => \N__13350\
        );

    \I__2929\ : ClkMux
    port map (
            O => \N__13535\,
            I => \N__13350\
        );

    \I__2928\ : ClkMux
    port map (
            O => \N__13534\,
            I => \N__13350\
        );

    \I__2927\ : ClkMux
    port map (
            O => \N__13533\,
            I => \N__13350\
        );

    \I__2926\ : ClkMux
    port map (
            O => \N__13532\,
            I => \N__13350\
        );

    \I__2925\ : ClkMux
    port map (
            O => \N__13531\,
            I => \N__13350\
        );

    \I__2924\ : ClkMux
    port map (
            O => \N__13530\,
            I => \N__13350\
        );

    \I__2923\ : ClkMux
    port map (
            O => \N__13529\,
            I => \N__13350\
        );

    \I__2922\ : ClkMux
    port map (
            O => \N__13528\,
            I => \N__13350\
        );

    \I__2921\ : ClkMux
    port map (
            O => \N__13527\,
            I => \N__13350\
        );

    \I__2920\ : ClkMux
    port map (
            O => \N__13526\,
            I => \N__13350\
        );

    \I__2919\ : ClkMux
    port map (
            O => \N__13525\,
            I => \N__13350\
        );

    \I__2918\ : ClkMux
    port map (
            O => \N__13524\,
            I => \N__13350\
        );

    \I__2917\ : ClkMux
    port map (
            O => \N__13523\,
            I => \N__13350\
        );

    \I__2916\ : ClkMux
    port map (
            O => \N__13522\,
            I => \N__13350\
        );

    \I__2915\ : ClkMux
    port map (
            O => \N__13521\,
            I => \N__13350\
        );

    \I__2914\ : ClkMux
    port map (
            O => \N__13520\,
            I => \N__13350\
        );

    \I__2913\ : ClkMux
    port map (
            O => \N__13519\,
            I => \N__13350\
        );

    \I__2912\ : ClkMux
    port map (
            O => \N__13518\,
            I => \N__13350\
        );

    \I__2911\ : ClkMux
    port map (
            O => \N__13517\,
            I => \N__13350\
        );

    \I__2910\ : ClkMux
    port map (
            O => \N__13516\,
            I => \N__13350\
        );

    \I__2909\ : ClkMux
    port map (
            O => \N__13515\,
            I => \N__13350\
        );

    \I__2908\ : ClkMux
    port map (
            O => \N__13514\,
            I => \N__13350\
        );

    \I__2907\ : ClkMux
    port map (
            O => \N__13513\,
            I => \N__13350\
        );

    \I__2906\ : ClkMux
    port map (
            O => \N__13512\,
            I => \N__13350\
        );

    \I__2905\ : ClkMux
    port map (
            O => \N__13511\,
            I => \N__13350\
        );

    \I__2904\ : ClkMux
    port map (
            O => \N__13510\,
            I => \N__13350\
        );

    \I__2903\ : ClkMux
    port map (
            O => \N__13509\,
            I => \N__13350\
        );

    \I__2902\ : ClkMux
    port map (
            O => \N__13508\,
            I => \N__13350\
        );

    \I__2901\ : ClkMux
    port map (
            O => \N__13507\,
            I => \N__13350\
        );

    \I__2900\ : ClkMux
    port map (
            O => \N__13506\,
            I => \N__13350\
        );

    \I__2899\ : ClkMux
    port map (
            O => \N__13505\,
            I => \N__13350\
        );

    \I__2898\ : ClkMux
    port map (
            O => \N__13504\,
            I => \N__13350\
        );

    \I__2897\ : ClkMux
    port map (
            O => \N__13503\,
            I => \N__13350\
        );

    \I__2896\ : ClkMux
    port map (
            O => \N__13502\,
            I => \N__13350\
        );

    \I__2895\ : ClkMux
    port map (
            O => \N__13501\,
            I => \N__13350\
        );

    \I__2894\ : ClkMux
    port map (
            O => \N__13500\,
            I => \N__13350\
        );

    \I__2893\ : ClkMux
    port map (
            O => \N__13499\,
            I => \N__13350\
        );

    \I__2892\ : ClkMux
    port map (
            O => \N__13498\,
            I => \N__13350\
        );

    \I__2891\ : ClkMux
    port map (
            O => \N__13497\,
            I => \N__13350\
        );

    \I__2890\ : ClkMux
    port map (
            O => \N__13496\,
            I => \N__13350\
        );

    \I__2889\ : ClkMux
    port map (
            O => \N__13495\,
            I => \N__13350\
        );

    \I__2888\ : ClkMux
    port map (
            O => \N__13494\,
            I => \N__13350\
        );

    \I__2887\ : ClkMux
    port map (
            O => \N__13493\,
            I => \N__13350\
        );

    \I__2886\ : ClkMux
    port map (
            O => \N__13492\,
            I => \N__13350\
        );

    \I__2885\ : ClkMux
    port map (
            O => \N__13491\,
            I => \N__13350\
        );

    \I__2884\ : ClkMux
    port map (
            O => \N__13490\,
            I => \N__13350\
        );

    \I__2883\ : ClkMux
    port map (
            O => \N__13489\,
            I => \N__13350\
        );

    \I__2882\ : ClkMux
    port map (
            O => \N__13488\,
            I => \N__13350\
        );

    \I__2881\ : ClkMux
    port map (
            O => \N__13487\,
            I => \N__13350\
        );

    \I__2880\ : ClkMux
    port map (
            O => \N__13486\,
            I => \N__13350\
        );

    \I__2879\ : ClkMux
    port map (
            O => \N__13485\,
            I => \N__13350\
        );

    \I__2878\ : ClkMux
    port map (
            O => \N__13484\,
            I => \N__13350\
        );

    \I__2877\ : ClkMux
    port map (
            O => \N__13483\,
            I => \N__13350\
        );

    \I__2876\ : GlobalMux
    port map (
            O => \N__13350\,
            I => \N__13347\
        );

    \I__2875\ : gio2CtrlBuf
    port map (
            O => \N__13347\,
            I => clk_g
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__13344\,
            I => \N__13341\
        );

    \I__2873\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13338\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__13338\,
            I => \N__13335\
        );

    \I__2871\ : Span12Mux_s4_h
    port map (
            O => \N__13335\,
            I => \N__13331\
        );

    \I__2870\ : InMux
    port map (
            O => \N__13334\,
            I => \N__13328\
        );

    \I__2869\ : Odrv12
    port map (
            O => \N__13331\,
            I => \Lab_UT.sec_clkD\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__13328\,
            I => \Lab_UT.sec_clkD\
        );

    \I__2867\ : InMux
    port map (
            O => \N__13323\,
            I => \N__13318\
        );

    \I__2866\ : InMux
    port map (
            O => \N__13322\,
            I => \N__13313\
        );

    \I__2865\ : InMux
    port map (
            O => \N__13321\,
            I => \N__13313\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__13318\,
            I => \N__13308\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__13313\,
            I => \N__13308\
        );

    \I__2862\ : Span4Mux_v
    port map (
            O => \N__13308\,
            I => \N__13303\
        );

    \I__2861\ : InMux
    port map (
            O => \N__13307\,
            I => \N__13298\
        );

    \I__2860\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13298\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__13303\,
            I => \Lab_UT.didpuu0.clkSecStrbZ0\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__13298\,
            I => \Lab_UT.didpuu0.clkSecStrbZ0\
        );

    \I__2857\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13290\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__13290\,
            I => \N__13287\
        );

    \I__2855\ : Span4Mux_h
    port map (
            O => \N__13287\,
            I => \N__13284\
        );

    \I__2854\ : Odrv4
    port map (
            O => \N__13284\,
            I => \L3_segment3_2\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__13281\,
            I => \L3_segment2_4_cascade_\
        );

    \I__2852\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13275\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__13275\,
            I => \N__13272\
        );

    \I__2850\ : Span4Mux_h
    port map (
            O => \N__13272\,
            I => \N__13269\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__13269\,
            I => \uu2.segment2_m_1Z0Z_6\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__13266\,
            I => \Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMUZ0Z_0_cascade_\
        );

    \I__2847\ : IoInMux
    port map (
            O => \N__13263\,
            I => \N__13260\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__13260\,
            I => \N__13257\
        );

    \I__2845\ : Span4Mux_s3_h
    port map (
            O => \N__13257\,
            I => \N__13254\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__13254\,
            I => led_c_3
        );

    \I__2843\ : InMux
    port map (
            O => \N__13251\,
            I => \N__13248\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__13248\,
            I => \Lab_UT.didpuu0.ledDisp00.selLed_RNI67CIZ0Z_0\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__13245\,
            I => \N__13241\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__13244\,
            I => \N__13238\
        );

    \I__2839\ : InMux
    port map (
            O => \N__13241\,
            I => \N__13233\
        );

    \I__2838\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13233\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__13233\,
            I => \N__13230\
        );

    \I__2836\ : Span4Mux_v
    port map (
            O => \N__13230\,
            I => \N__13226\
        );

    \I__2835\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13223\
        );

    \I__2834\ : Odrv4
    port map (
            O => \N__13226\,
            I => \Lab_UT.un11_segmentUQ_1\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__13223\,
            I => \Lab_UT.un11_segmentUQ_1\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__13218\,
            I => \Lab_UT.didpuu0.countEnMtens_0_a4_0_cascade_\
        );

    \I__2831\ : InMux
    port map (
            O => \N__13215\,
            I => \N__13211\
        );

    \I__2830\ : InMux
    port map (
            O => \N__13214\,
            I => \N__13208\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__13211\,
            I => \N__13205\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__13208\,
            I => \N__13202\
        );

    \I__2827\ : Span4Mux_v
    port map (
            O => \N__13205\,
            I => \N__13199\
        );

    \I__2826\ : Span4Mux_v
    port map (
            O => \N__13202\,
            I => \N__13194\
        );

    \I__2825\ : Span4Mux_h
    port map (
            O => \N__13199\,
            I => \N__13194\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__13194\,
            I => \Lab_UT.didpuu0.countEnMtens_0_a4_1\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__13191\,
            I => \Lab_UT.didpuu0.countEnMtens_0_a4_1_cascade_\
        );

    \I__2822\ : InMux
    port map (
            O => \N__13188\,
            I => \N__13185\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__13185\,
            I => \N__13180\
        );

    \I__2820\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13174\
        );

    \I__2819\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13171\
        );

    \I__2818\ : Span4Mux_v
    port map (
            O => \N__13180\,
            I => \N__13168\
        );

    \I__2817\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13161\
        );

    \I__2816\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13161\
        );

    \I__2815\ : InMux
    port map (
            O => \N__13177\,
            I => \N__13161\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__13174\,
            I => \Lab_UT.didpuu0.countEnStens\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__13171\,
            I => \Lab_UT.didpuu0.countEnStens\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__13168\,
            I => \Lab_UT.didpuu0.countEnStens\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__13161\,
            I => \Lab_UT.didpuu0.countEnStens\
        );

    \I__2810\ : InMux
    port map (
            O => \N__13152\,
            I => \N__13148\
        );

    \I__2809\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13145\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__13148\,
            I => \N__13142\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__13145\,
            I => \N__13139\
        );

    \I__2806\ : Span4Mux_h
    port map (
            O => \N__13142\,
            I => \N__13136\
        );

    \I__2805\ : Sp12to4
    port map (
            O => \N__13139\,
            I => \N__13133\
        );

    \I__2804\ : Span4Mux_v
    port map (
            O => \N__13136\,
            I => \N__13130\
        );

    \I__2803\ : Odrv12
    port map (
            O => \N__13133\,
            I => \Lab_UT.didpuu0.countEnMtens\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__13130\,
            I => \Lab_UT.didpuu0.countEnMtens\
        );

    \I__2801\ : InMux
    port map (
            O => \N__13125\,
            I => \N__13122\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__13122\,
            I => \Lab_UT.un152_segmentUQ_1\
        );

    \I__2799\ : CEMux
    port map (
            O => \N__13119\,
            I => \N__13116\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__13116\,
            I => \N__13113\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__13113\,
            I => \N__13110\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__13110\,
            I => \Lab_UT.didpuu0.didpstens.countEnStens_0\
        );

    \I__2795\ : InMux
    port map (
            O => \N__13107\,
            I => \N__13104\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__13104\,
            I => \uu2.un1_segment4_3_bmZ0\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__13101\,
            I => \uu2.un1_segment4_3_amZ0_cascade_\
        );

    \I__2792\ : InMux
    port map (
            O => \N__13098\,
            I => \N__13095\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__13095\,
            I => \uu2.un1_segment4_9_ns_1\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__13092\,
            I => \uu2.N_289_cascade_\
        );

    \I__2789\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13086\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__13086\,
            I => \uu2.w_addr_displaying_fast_RNIFU9M8Z0Z_8\
        );

    \I__2787\ : InMux
    port map (
            O => \N__13083\,
            I => \N__13078\
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__13082\,
            I => \N__13074\
        );

    \I__2785\ : InMux
    port map (
            O => \N__13081\,
            I => \N__13071\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__13078\,
            I => \N__13066\
        );

    \I__2783\ : InMux
    port map (
            O => \N__13077\,
            I => \N__13061\
        );

    \I__2782\ : InMux
    port map (
            O => \N__13074\,
            I => \N__13061\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__13071\,
            I => \N__13057\
        );

    \I__2780\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13052\
        );

    \I__2779\ : InMux
    port map (
            O => \N__13069\,
            I => \N__13052\
        );

    \I__2778\ : Span4Mux_h
    port map (
            O => \N__13066\,
            I => \N__13047\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__13061\,
            I => \N__13047\
        );

    \I__2776\ : InMux
    port map (
            O => \N__13060\,
            I => \N__13044\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__13057\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__13052\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__13047\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__13044\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__13035\,
            I => \N__13032\
        );

    \I__2770\ : InMux
    port map (
            O => \N__13032\,
            I => \N__13029\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__13029\,
            I => \N__13026\
        );

    \I__2768\ : Span4Mux_h
    port map (
            O => \N__13026\,
            I => \N__13023\
        );

    \I__2767\ : Odrv4
    port map (
            O => \N__13023\,
            I => \uu2.N_1\
        );

    \I__2766\ : InMux
    port map (
            O => \N__13020\,
            I => \N__13017\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__13017\,
            I => \uu2.w_addr_displaying_4_rep1_RNIAVDBZ0Z_0\
        );

    \I__2764\ : InMux
    port map (
            O => \N__13014\,
            I => \N__13011\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__13011\,
            I => \N__13008\
        );

    \I__2762\ : Span4Mux_h
    port map (
            O => \N__13008\,
            I => \N__13005\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__13005\,
            I => \uu2.w_addr_displaying_fast_RNIKFIEZ0Z_6\
        );

    \I__2760\ : InMux
    port map (
            O => \N__13002\,
            I => \N__12999\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__12999\,
            I => \N__12996\
        );

    \I__2758\ : Span4Mux_h
    port map (
            O => \N__12996\,
            I => \N__12993\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__12993\,
            I => \uu2.w_addr_displaying_fast_RNIN0TSZ0Z_4\
        );

    \I__2756\ : InMux
    port map (
            O => \N__12990\,
            I => \N__12980\
        );

    \I__2755\ : InMux
    port map (
            O => \N__12989\,
            I => \N__12980\
        );

    \I__2754\ : InMux
    port map (
            O => \N__12988\,
            I => \N__12977\
        );

    \I__2753\ : InMux
    port map (
            O => \N__12987\,
            I => \N__12970\
        );

    \I__2752\ : InMux
    port map (
            O => \N__12986\,
            I => \N__12970\
        );

    \I__2751\ : InMux
    port map (
            O => \N__12985\,
            I => \N__12970\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__12980\,
            I => \uu2.w_addr_displaying_fastZ0Z_4\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__12977\,
            I => \uu2.w_addr_displaying_fastZ0Z_4\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__12970\,
            I => \uu2.w_addr_displaying_fastZ0Z_4\
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__12963\,
            I => \N__12958\
        );

    \I__2746\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12955\
        );

    \I__2745\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12949\
        );

    \I__2744\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12946\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__12955\,
            I => \N__12943\
        );

    \I__2742\ : InMux
    port map (
            O => \N__12954\,
            I => \N__12940\
        );

    \I__2741\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12935\
        );

    \I__2740\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12935\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__12949\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__12946\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__12943\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__12940\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__12935\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2734\ : InMux
    port map (
            O => \N__12924\,
            I => \N__12921\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__12921\,
            I => \uu2.N_10_0\
        );

    \I__2732\ : CascadeMux
    port map (
            O => \N__12918\,
            I => \N__12914\
        );

    \I__2731\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12911\
        );

    \I__2730\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12908\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__12911\,
            I => \N__12905\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__12908\,
            I => \N__12902\
        );

    \I__2727\ : Span4Mux_h
    port map (
            O => \N__12905\,
            I => \N__12899\
        );

    \I__2726\ : Span4Mux_h
    port map (
            O => \N__12902\,
            I => \N__12894\
        );

    \I__2725\ : Span4Mux_v
    port map (
            O => \N__12899\,
            I => \N__12894\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__12894\,
            I => \Lab_UT.didpuu0.didpsones.N_38\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__12891\,
            I => \N__12888\
        );

    \I__2722\ : InMux
    port map (
            O => \N__12888\,
            I => \N__12885\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__12885\,
            I => \N__12882\
        );

    \I__2720\ : Span4Mux_v
    port map (
            O => \N__12882\,
            I => \N__12879\
        );

    \I__2719\ : Span4Mux_s3_h
    port map (
            O => \N__12879\,
            I => \N__12876\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__12876\,
            I => \Lab_UT.didpuu0.didpsones.N_32\
        );

    \I__2717\ : InMux
    port map (
            O => \N__12873\,
            I => \N__12869\
        );

    \I__2716\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12865\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__12869\,
            I => \N__12862\
        );

    \I__2714\ : InMux
    port map (
            O => \N__12868\,
            I => \N__12859\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__12865\,
            I => \N__12856\
        );

    \I__2712\ : Span4Mux_h
    port map (
            O => \N__12862\,
            I => \N__12849\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__12859\,
            I => \N__12849\
        );

    \I__2710\ : Span4Mux_h
    port map (
            O => \N__12856\,
            I => \N__12849\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__12849\,
            I => \Lab_UT_dec0_un137_segmentUQ\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__12846\,
            I => \uu2.segment1_m_2Z0Z_0_cascade_\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__12843\,
            I => \uu2.segment1_m_0_cascade_\
        );

    \I__2706\ : InMux
    port map (
            O => \N__12840\,
            I => \N__12831\
        );

    \I__2705\ : InMux
    port map (
            O => \N__12839\,
            I => \N__12826\
        );

    \I__2704\ : InMux
    port map (
            O => \N__12838\,
            I => \N__12826\
        );

    \I__2703\ : InMux
    port map (
            O => \N__12837\,
            I => \N__12823\
        );

    \I__2702\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12820\
        );

    \I__2701\ : InMux
    port map (
            O => \N__12835\,
            I => \N__12814\
        );

    \I__2700\ : InMux
    port map (
            O => \N__12834\,
            I => \N__12814\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__12831\,
            I => \N__12805\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__12826\,
            I => \N__12805\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__12823\,
            I => \N__12800\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__12820\,
            I => \N__12800\
        );

    \I__2695\ : InMux
    port map (
            O => \N__12819\,
            I => \N__12791\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__12814\,
            I => \N__12788\
        );

    \I__2693\ : InMux
    port map (
            O => \N__12813\,
            I => \N__12779\
        );

    \I__2692\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12779\
        );

    \I__2691\ : InMux
    port map (
            O => \N__12811\,
            I => \N__12779\
        );

    \I__2690\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12779\
        );

    \I__2689\ : Span4Mux_v
    port map (
            O => \N__12805\,
            I => \N__12774\
        );

    \I__2688\ : Span4Mux_h
    port map (
            O => \N__12800\,
            I => \N__12774\
        );

    \I__2687\ : InMux
    port map (
            O => \N__12799\,
            I => \N__12767\
        );

    \I__2686\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12767\
        );

    \I__2685\ : InMux
    port map (
            O => \N__12797\,
            I => \N__12767\
        );

    \I__2684\ : InMux
    port map (
            O => \N__12796\,
            I => \N__12764\
        );

    \I__2683\ : InMux
    port map (
            O => \N__12795\,
            I => \N__12761\
        );

    \I__2682\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12758\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__12791\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__12788\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__12779\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__12774\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__12767\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__12764\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__12761\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__12758\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2673\ : InMux
    port map (
            O => \N__12741\,
            I => \N__12738\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__12738\,
            I => \uu2.segment3_m_6\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__12735\,
            I => \uu2.un1_segment1_iv_0_cascade_\
        );

    \I__2670\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12724\
        );

    \I__2669\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12719\
        );

    \I__2668\ : InMux
    port map (
            O => \N__12730\,
            I => \N__12719\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__12729\,
            I => \N__12716\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__12728\,
            I => \N__12712\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__12727\,
            I => \N__12709\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__12724\,
            I => \N__12704\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__12719\,
            I => \N__12704\
        );

    \I__2662\ : InMux
    port map (
            O => \N__12716\,
            I => \N__12699\
        );

    \I__2661\ : InMux
    port map (
            O => \N__12715\,
            I => \N__12699\
        );

    \I__2660\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12694\
        );

    \I__2659\ : InMux
    port map (
            O => \N__12709\,
            I => \N__12694\
        );

    \I__2658\ : Span4Mux_h
    port map (
            O => \N__12704\,
            I => \N__12691\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__12699\,
            I => \N__12686\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__12694\,
            I => \N__12686\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__12691\,
            I => \uu2.un1_segment1_0\
        );

    \I__2654\ : Odrv4
    port map (
            O => \N__12686\,
            I => \uu2.un1_segment1_0\
        );

    \I__2653\ : InMux
    port map (
            O => \N__12681\,
            I => \N__12678\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__12678\,
            I => \uu2.un1_segment4_sn_N_61\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__12675\,
            I => \uu2.w_addr_displaying_fast_RNI6N2KZ0Z_5_cascade_\
        );

    \I__2650\ : InMux
    port map (
            O => \N__12672\,
            I => \N__12669\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__12669\,
            I => \uu2.w_addr_displaying_fast_RNID5QHZ0Z_5\
        );

    \I__2648\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12663\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__12663\,
            I => \N__12660\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__12660\,
            I => \uu2.un1_segment4_sn_N_39_0\
        );

    \I__2645\ : InMux
    port map (
            O => \N__12657\,
            I => \N__12654\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__12654\,
            I => \N__12651\
        );

    \I__2643\ : Odrv12
    port map (
            O => \N__12651\,
            I => \uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__12648\,
            I => \uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4_cascade_\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__12645\,
            I => \N__12640\
        );

    \I__2640\ : InMux
    port map (
            O => \N__12644\,
            I => \N__12635\
        );

    \I__2639\ : InMux
    port map (
            O => \N__12643\,
            I => \N__12635\
        );

    \I__2638\ : InMux
    port map (
            O => \N__12640\,
            I => \N__12632\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__12635\,
            I => \N__12627\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__12632\,
            I => \N__12624\
        );

    \I__2635\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12619\
        );

    \I__2634\ : InMux
    port map (
            O => \N__12630\,
            I => \N__12619\
        );

    \I__2633\ : Span4Mux_h
    port map (
            O => \N__12627\,
            I => \N__12614\
        );

    \I__2632\ : Span4Mux_h
    port map (
            O => \N__12624\,
            I => \N__12609\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__12619\,
            I => \N__12609\
        );

    \I__2630\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12604\
        );

    \I__2629\ : InMux
    port map (
            O => \N__12617\,
            I => \N__12604\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__12614\,
            I => \uu2.w_addr_displaying_RNILB202Z0Z_4\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__12609\,
            I => \uu2.w_addr_displaying_RNILB202Z0Z_4\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__12604\,
            I => \uu2.w_addr_displaying_RNILB202Z0Z_4\
        );

    \I__2625\ : InMux
    port map (
            O => \N__12597\,
            I => \N__12594\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__12594\,
            I => \N__12591\
        );

    \I__2623\ : Span4Mux_h
    port map (
            O => \N__12591\,
            I => \N__12588\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__12588\,
            I => \uu2.N_92\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__12585\,
            I => \N__12582\
        );

    \I__2620\ : InMux
    port map (
            O => \N__12582\,
            I => \N__12579\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__12579\,
            I => \uu2.w_addr_displaying_4_0_i_fast_6\
        );

    \I__2618\ : InMux
    port map (
            O => \N__12576\,
            I => \N__12572\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__12575\,
            I => \N__12566\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__12572\,
            I => \N__12558\
        );

    \I__2615\ : InMux
    port map (
            O => \N__12571\,
            I => \N__12551\
        );

    \I__2614\ : InMux
    port map (
            O => \N__12570\,
            I => \N__12551\
        );

    \I__2613\ : InMux
    port map (
            O => \N__12569\,
            I => \N__12551\
        );

    \I__2612\ : InMux
    port map (
            O => \N__12566\,
            I => \N__12548\
        );

    \I__2611\ : InMux
    port map (
            O => \N__12565\,
            I => \N__12545\
        );

    \I__2610\ : InMux
    port map (
            O => \N__12564\,
            I => \N__12540\
        );

    \I__2609\ : InMux
    port map (
            O => \N__12563\,
            I => \N__12540\
        );

    \I__2608\ : InMux
    port map (
            O => \N__12562\,
            I => \N__12535\
        );

    \I__2607\ : InMux
    port map (
            O => \N__12561\,
            I => \N__12535\
        );

    \I__2606\ : Span4Mux_h
    port map (
            O => \N__12558\,
            I => \N__12531\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__12551\,
            I => \N__12528\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__12548\,
            I => \N__12525\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__12545\,
            I => \N__12516\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__12540\,
            I => \N__12516\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__12535\,
            I => \N__12516\
        );

    \I__2600\ : InMux
    port map (
            O => \N__12534\,
            I => \N__12513\
        );

    \I__2599\ : Span4Mux_h
    port map (
            O => \N__12531\,
            I => \N__12510\
        );

    \I__2598\ : Span4Mux_v
    port map (
            O => \N__12528\,
            I => \N__12505\
        );

    \I__2597\ : Span4Mux_h
    port map (
            O => \N__12525\,
            I => \N__12505\
        );

    \I__2596\ : InMux
    port map (
            O => \N__12524\,
            I => \N__12500\
        );

    \I__2595\ : InMux
    port map (
            O => \N__12523\,
            I => \N__12500\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__12516\,
            I => \N__12497\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__12513\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__12510\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__12505\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__12500\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__12497\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__12486\,
            I => \uu2.un15_w_data_displaying_cascade_\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__12483\,
            I => \N__12479\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__12482\,
            I => \N__12472\
        );

    \I__2585\ : InMux
    port map (
            O => \N__12479\,
            I => \N__12463\
        );

    \I__2584\ : InMux
    port map (
            O => \N__12478\,
            I => \N__12451\
        );

    \I__2583\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12451\
        );

    \I__2582\ : InMux
    port map (
            O => \N__12476\,
            I => \N__12451\
        );

    \I__2581\ : InMux
    port map (
            O => \N__12475\,
            I => \N__12451\
        );

    \I__2580\ : InMux
    port map (
            O => \N__12472\,
            I => \N__12448\
        );

    \I__2579\ : InMux
    port map (
            O => \N__12471\,
            I => \N__12445\
        );

    \I__2578\ : InMux
    port map (
            O => \N__12470\,
            I => \N__12440\
        );

    \I__2577\ : InMux
    port map (
            O => \N__12469\,
            I => \N__12440\
        );

    \I__2576\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12433\
        );

    \I__2575\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12433\
        );

    \I__2574\ : InMux
    port map (
            O => \N__12466\,
            I => \N__12433\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__12463\,
            I => \N__12430\
        );

    \I__2572\ : CascadeMux
    port map (
            O => \N__12462\,
            I => \N__12421\
        );

    \I__2571\ : InMux
    port map (
            O => \N__12461\,
            I => \N__12415\
        );

    \I__2570\ : InMux
    port map (
            O => \N__12460\,
            I => \N__12415\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__12451\,
            I => \N__12412\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__12448\,
            I => \N__12405\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__12445\,
            I => \N__12405\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__12440\,
            I => \N__12405\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__12433\,
            I => \N__12400\
        );

    \I__2564\ : Span4Mux_v
    port map (
            O => \N__12430\,
            I => \N__12400\
        );

    \I__2563\ : InMux
    port map (
            O => \N__12429\,
            I => \N__12392\
        );

    \I__2562\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12392\
        );

    \I__2561\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12392\
        );

    \I__2560\ : InMux
    port map (
            O => \N__12426\,
            I => \N__12389\
        );

    \I__2559\ : InMux
    port map (
            O => \N__12425\,
            I => \N__12386\
        );

    \I__2558\ : InMux
    port map (
            O => \N__12424\,
            I => \N__12379\
        );

    \I__2557\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12379\
        );

    \I__2556\ : InMux
    port map (
            O => \N__12420\,
            I => \N__12379\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__12415\,
            I => \N__12376\
        );

    \I__2554\ : Span4Mux_v
    port map (
            O => \N__12412\,
            I => \N__12371\
        );

    \I__2553\ : Span4Mux_v
    port map (
            O => \N__12405\,
            I => \N__12371\
        );

    \I__2552\ : Span4Mux_h
    port map (
            O => \N__12400\,
            I => \N__12368\
        );

    \I__2551\ : InMux
    port map (
            O => \N__12399\,
            I => \N__12365\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__12392\,
            I => \N__12360\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__12389\,
            I => \N__12360\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__12386\,
            I => \uu2.un19_w_addr_userZ0Z_0\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__12379\,
            I => \uu2.un19_w_addr_userZ0Z_0\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__12376\,
            I => \uu2.un19_w_addr_userZ0Z_0\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__12371\,
            I => \uu2.un19_w_addr_userZ0Z_0\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__12368\,
            I => \uu2.un19_w_addr_userZ0Z_0\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__12365\,
            I => \uu2.un19_w_addr_userZ0Z_0\
        );

    \I__2542\ : Odrv12
    port map (
            O => \N__12360\,
            I => \uu2.un19_w_addr_userZ0Z_0\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__12345\,
            I => \uu2.un21_w_addr_displaying_i_cascade_\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__12342\,
            I => \N__12339\
        );

    \I__2539\ : InMux
    port map (
            O => \N__12339\,
            I => \N__12334\
        );

    \I__2538\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12329\
        );

    \I__2537\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12329\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__12334\,
            I => \uu2.un15_w_data_displaying\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__12329\,
            I => \uu2.un15_w_data_displaying\
        );

    \I__2534\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12317\
        );

    \I__2533\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12317\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__12322\,
            I => \N__12312\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__12317\,
            I => \N__12309\
        );

    \I__2530\ : InMux
    port map (
            O => \N__12316\,
            I => \N__12306\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__12315\,
            I => \N__12302\
        );

    \I__2528\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12299\
        );

    \I__2527\ : Span4Mux_h
    port map (
            O => \N__12309\,
            I => \N__12294\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__12306\,
            I => \N__12294\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__12305\,
            I => \N__12288\
        );

    \I__2524\ : InMux
    port map (
            O => \N__12302\,
            I => \N__12285\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__12299\,
            I => \N__12282\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__12294\,
            I => \N__12279\
        );

    \I__2521\ : InMux
    port map (
            O => \N__12293\,
            I => \N__12276\
        );

    \I__2520\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12269\
        );

    \I__2519\ : InMux
    port map (
            O => \N__12291\,
            I => \N__12269\
        );

    \I__2518\ : InMux
    port map (
            O => \N__12288\,
            I => \N__12269\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__12285\,
            I => \N__12266\
        );

    \I__2516\ : Span4Mux_h
    port map (
            O => \N__12282\,
            I => \N__12263\
        );

    \I__2515\ : Odrv4
    port map (
            O => \N__12279\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__12276\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__12269\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2512\ : Odrv12
    port map (
            O => \N__12266\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2511\ : Odrv4
    port map (
            O => \N__12263\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2510\ : InMux
    port map (
            O => \N__12252\,
            I => \N__12249\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__12249\,
            I => \uu2.w_addr_displaying_4_0_i_rep1_6\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__12246\,
            I => \uu2.w_addr_displaying_5_rep1_RNI3HMTZ0_cascade_\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__12243\,
            I => \Lab_UT.didpuu0.countEnStens_cascade_\
        );

    \I__2506\ : InMux
    port map (
            O => \N__12240\,
            I => \N__12237\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__12237\,
            I => \uu2.un1_segment4_2_amZ0Z_1\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__12234\,
            I => \uu2.w_addr_displaying_4_0_i_6_cascade_\
        );

    \I__2503\ : InMux
    port map (
            O => \N__12231\,
            I => \N__12226\
        );

    \I__2502\ : InMux
    port map (
            O => \N__12230\,
            I => \N__12217\
        );

    \I__2501\ : InMux
    port map (
            O => \N__12229\,
            I => \N__12217\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__12226\,
            I => \N__12214\
        );

    \I__2499\ : CascadeMux
    port map (
            O => \N__12225\,
            I => \N__12209\
        );

    \I__2498\ : InMux
    port map (
            O => \N__12224\,
            I => \N__12204\
        );

    \I__2497\ : InMux
    port map (
            O => \N__12223\,
            I => \N__12204\
        );

    \I__2496\ : InMux
    port map (
            O => \N__12222\,
            I => \N__12201\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__12217\,
            I => \N__12198\
        );

    \I__2494\ : Span4Mux_v
    port map (
            O => \N__12214\,
            I => \N__12195\
        );

    \I__2493\ : InMux
    port map (
            O => \N__12213\,
            I => \N__12192\
        );

    \I__2492\ : InMux
    port map (
            O => \N__12212\,
            I => \N__12187\
        );

    \I__2491\ : InMux
    port map (
            O => \N__12209\,
            I => \N__12187\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__12204\,
            I => \N__12182\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__12201\,
            I => \N__12182\
        );

    \I__2488\ : Span4Mux_h
    port map (
            O => \N__12198\,
            I => \N__12178\
        );

    \I__2487\ : Span4Mux_h
    port map (
            O => \N__12195\,
            I => \N__12173\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__12192\,
            I => \N__12173\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__12187\,
            I => \N__12168\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__12182\,
            I => \N__12168\
        );

    \I__2483\ : InMux
    port map (
            O => \N__12181\,
            I => \N__12165\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__12178\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__12173\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__12168\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__12165\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__12156\,
            I => \N__12153\
        );

    \I__2477\ : InMux
    port map (
            O => \N__12153\,
            I => \N__12150\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__12150\,
            I => \N__12147\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__12147\,
            I => \uu2.g0_i_o4_0_a8_3_1\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__12144\,
            I => \uu2_un3_r_clk_en_0_cascade_\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__12141\,
            I => \N__12138\
        );

    \I__2472\ : InMux
    port map (
            O => \N__12138\,
            I => \N__12135\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__12135\,
            I => \uu2.un349_ci_0\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__12132\,
            I => \N__12127\
        );

    \I__2469\ : InMux
    port map (
            O => \N__12131\,
            I => \N__12124\
        );

    \I__2468\ : InMux
    port map (
            O => \N__12130\,
            I => \N__12119\
        );

    \I__2467\ : InMux
    port map (
            O => \N__12127\,
            I => \N__12119\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__12124\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__12119\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__2464\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12105\
        );

    \I__2463\ : InMux
    port map (
            O => \N__12113\,
            I => \N__12105\
        );

    \I__2462\ : InMux
    port map (
            O => \N__12112\,
            I => \N__12105\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__12105\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__12102\,
            I => \N__12098\
        );

    \I__2459\ : InMux
    port map (
            O => \N__12101\,
            I => \N__12094\
        );

    \I__2458\ : InMux
    port map (
            O => \N__12098\,
            I => \N__12089\
        );

    \I__2457\ : InMux
    port map (
            O => \N__12097\,
            I => \N__12089\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__12094\,
            I => \N__12086\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__12089\,
            I => \N__12083\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__12086\,
            I => \uu2.vbuf_count.un382_ci_8_1\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__12083\,
            I => \uu2.vbuf_count.un382_ci_8_1\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__12078\,
            I => \N__12072\
        );

    \I__2451\ : InMux
    port map (
            O => \N__12077\,
            I => \N__12069\
        );

    \I__2450\ : InMux
    port map (
            O => \N__12076\,
            I => \N__12064\
        );

    \I__2449\ : InMux
    port map (
            O => \N__12075\,
            I => \N__12064\
        );

    \I__2448\ : InMux
    port map (
            O => \N__12072\,
            I => \N__12061\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__12069\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__12064\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__12061\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__12054\,
            I => \N__12049\
        );

    \I__2443\ : InMux
    port map (
            O => \N__12053\,
            I => \N__12041\
        );

    \I__2442\ : InMux
    port map (
            O => \N__12052\,
            I => \N__12041\
        );

    \I__2441\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12041\
        );

    \I__2440\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12036\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__12041\,
            I => \N__12033\
        );

    \I__2438\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12028\
        );

    \I__2437\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12028\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__12036\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__12033\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__12028\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__12021\,
            I => \N__12018\
        );

    \I__2432\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12013\
        );

    \I__2431\ : InMux
    port map (
            O => \N__12017\,
            I => \N__12010\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__12016\,
            I => \N__12003\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__12013\,
            I => \N__11998\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__12010\,
            I => \N__11998\
        );

    \I__2427\ : InMux
    port map (
            O => \N__12009\,
            I => \N__11995\
        );

    \I__2426\ : InMux
    port map (
            O => \N__12008\,
            I => \N__11986\
        );

    \I__2425\ : InMux
    port map (
            O => \N__12007\,
            I => \N__11986\
        );

    \I__2424\ : InMux
    port map (
            O => \N__12006\,
            I => \N__11986\
        );

    \I__2423\ : InMux
    port map (
            O => \N__12003\,
            I => \N__11986\
        );

    \I__2422\ : Odrv4
    port map (
            O => \N__11998\,
            I => \uu2.un316_ci\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__11995\,
            I => \uu2.un316_ci\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__11986\,
            I => \uu2.un316_ci\
        );

    \I__2419\ : InMux
    port map (
            O => \N__11979\,
            I => \N__11972\
        );

    \I__2418\ : InMux
    port map (
            O => \N__11978\,
            I => \N__11967\
        );

    \I__2417\ : InMux
    port map (
            O => \N__11977\,
            I => \N__11967\
        );

    \I__2416\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11962\
        );

    \I__2415\ : InMux
    port map (
            O => \N__11975\,
            I => \N__11962\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__11972\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__11967\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__11962\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__2411\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11949\
        );

    \I__2410\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11946\
        );

    \I__2409\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11943\
        );

    \I__2408\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11940\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__11949\,
            I => \N__11937\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__11946\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__11943\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__11940\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__11937\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__2402\ : InMux
    port map (
            O => \N__11928\,
            I => \N__11925\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__11925\,
            I => \uu2.un382_ci\
        );

    \I__2400\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11915\
        );

    \I__2399\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11910\
        );

    \I__2398\ : InMux
    port map (
            O => \N__11920\,
            I => \N__11907\
        );

    \I__2397\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11904\
        );

    \I__2396\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11901\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__11915\,
            I => \N__11898\
        );

    \I__2394\ : InMux
    port map (
            O => \N__11914\,
            I => \N__11893\
        );

    \I__2393\ : InMux
    port map (
            O => \N__11913\,
            I => \N__11893\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__11910\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__11907\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__11904\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__11901\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__11898\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__11893\,
            I => uu2_un3_r_clk_en_0
        );

    \I__2386\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11876\
        );

    \I__2385\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11873\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__11876\,
            I => \uu2.l_countZ0Z_10\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__11873\,
            I => \uu2.l_countZ0Z_10\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__11868\,
            I => \Lab_UT.didpuu0.countEnMones_cascade_\
        );

    \I__2381\ : CEMux
    port map (
            O => \N__11865\,
            I => \N__11862\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__11862\,
            I => \N__11859\
        );

    \I__2379\ : Span4Mux_h
    port map (
            O => \N__11859\,
            I => \N__11856\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__11856\,
            I => \N__11853\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__11853\,
            I => \Lab_UT.didpuu0.didpmones.countEnMones_0\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__11850\,
            I => \N__11845\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__11849\,
            I => \N__11842\
        );

    \I__2374\ : InMux
    port map (
            O => \N__11848\,
            I => \N__11836\
        );

    \I__2373\ : InMux
    port map (
            O => \N__11845\,
            I => \N__11836\
        );

    \I__2372\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11831\
        );

    \I__2371\ : InMux
    port map (
            O => \N__11841\,
            I => \N__11831\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__11836\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__11831\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__2368\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11812\
        );

    \I__2367\ : InMux
    port map (
            O => \N__11825\,
            I => \N__11812\
        );

    \I__2366\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11812\
        );

    \I__2365\ : InMux
    port map (
            O => \N__11823\,
            I => \N__11812\
        );

    \I__2364\ : InMux
    port map (
            O => \N__11822\,
            I => \N__11807\
        );

    \I__2363\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11807\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__11812\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__11807\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__11802\,
            I => \N__11799\
        );

    \I__2359\ : InMux
    port map (
            O => \N__11799\,
            I => \N__11792\
        );

    \I__2358\ : InMux
    port map (
            O => \N__11798\,
            I => \N__11792\
        );

    \I__2357\ : InMux
    port map (
            O => \N__11797\,
            I => \N__11789\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__11792\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__11789\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__2354\ : InMux
    port map (
            O => \N__11784\,
            I => \N__11771\
        );

    \I__2353\ : InMux
    port map (
            O => \N__11783\,
            I => \N__11771\
        );

    \I__2352\ : InMux
    port map (
            O => \N__11782\,
            I => \N__11771\
        );

    \I__2351\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11771\
        );

    \I__2350\ : InMux
    port map (
            O => \N__11780\,
            I => \N__11768\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__11771\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__11768\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__2347\ : InMux
    port map (
            O => \N__11763\,
            I => \N__11760\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__11760\,
            I => \uu2.un3_r_clk_en_7\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__11757\,
            I => \uu2.un3_r_clk_en_0_0_cascade_\
        );

    \I__2344\ : InMux
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__11751\,
            I => \uu2.un3_r_clk_en_6\
        );

    \I__2342\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11745\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__11745\,
            I => \N__11742\
        );

    \I__2340\ : Span12Mux_s6_h
    port map (
            O => \N__11742\,
            I => \N__11739\
        );

    \I__2339\ : Odrv12
    port map (
            O => \N__11739\,
            I => \uu2.mem0.G_14_0_a6_2_1\
        );

    \I__2338\ : InMux
    port map (
            O => \N__11736\,
            I => \N__11733\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__11733\,
            I => \uu2.mem0.bitmap_pmux_1_1_2_tz_0\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__11730\,
            I => \N__11727\
        );

    \I__2335\ : InMux
    port map (
            O => \N__11727\,
            I => \N__11724\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__11724\,
            I => \uu2.bitmap_pmux_1_1_2_tz_1_0\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__11721\,
            I => \uu2.bitmap_pmux_1_1_2_tz_1_0_cascade_\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__11718\,
            I => \uu2.mem0.bitmap_pmux_1_1_2_tz_cascade_\
        );

    \I__2331\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11712\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__11712\,
            I => \N__11709\
        );

    \I__2329\ : Span4Mux_v
    port map (
            O => \N__11709\,
            I => \N__11706\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__11706\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_33\
        );

    \I__2327\ : InMux
    port map (
            O => \N__11703\,
            I => \N__11700\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__11700\,
            I => \N__11695\
        );

    \I__2325\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11691\
        );

    \I__2324\ : InMux
    port map (
            O => \N__11698\,
            I => \N__11688\
        );

    \I__2323\ : Span4Mux_h
    port map (
            O => \N__11695\,
            I => \N__11680\
        );

    \I__2322\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11677\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__11691\,
            I => \N__11674\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__11688\,
            I => \N__11671\
        );

    \I__2319\ : InMux
    port map (
            O => \N__11687\,
            I => \N__11664\
        );

    \I__2318\ : InMux
    port map (
            O => \N__11686\,
            I => \N__11664\
        );

    \I__2317\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11664\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__11684\,
            I => \N__11658\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__11683\,
            I => \N__11655\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__11680\,
            I => \N__11652\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__11677\,
            I => \N__11649\
        );

    \I__2312\ : Span4Mux_v
    port map (
            O => \N__11674\,
            I => \N__11642\
        );

    \I__2311\ : Span4Mux_h
    port map (
            O => \N__11671\,
            I => \N__11642\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__11664\,
            I => \N__11642\
        );

    \I__2309\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11631\
        );

    \I__2308\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11631\
        );

    \I__2307\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11631\
        );

    \I__2306\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11631\
        );

    \I__2305\ : InMux
    port map (
            O => \N__11655\,
            I => \N__11631\
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__11652\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2303\ : Odrv4
    port map (
            O => \N__11649\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__11642\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__11631\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__11622\,
            I => \uu2.w_addr_displaying_RNI8NHB1Z0Z_2_cascade_\
        );

    \I__2299\ : InMux
    port map (
            O => \N__11619\,
            I => \N__11616\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__11616\,
            I => \N__11613\
        );

    \I__2297\ : Span4Mux_v
    port map (
            O => \N__11613\,
            I => \N__11610\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__11610\,
            I => \uu2.w_addr_displaying_RNI18582Z0Z_8\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__11607\,
            I => \N__11603\
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__11606\,
            I => \N__11600\
        );

    \I__2293\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11590\
        );

    \I__2292\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11590\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__11599\,
            I => \N__11583\
        );

    \I__2290\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11580\
        );

    \I__2289\ : InMux
    port map (
            O => \N__11597\,
            I => \N__11575\
        );

    \I__2288\ : InMux
    port map (
            O => \N__11596\,
            I => \N__11575\
        );

    \I__2287\ : InMux
    port map (
            O => \N__11595\,
            I => \N__11572\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__11590\,
            I => \N__11569\
        );

    \I__2285\ : InMux
    port map (
            O => \N__11589\,
            I => \N__11562\
        );

    \I__2284\ : InMux
    port map (
            O => \N__11588\,
            I => \N__11562\
        );

    \I__2283\ : InMux
    port map (
            O => \N__11587\,
            I => \N__11562\
        );

    \I__2282\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11557\
        );

    \I__2281\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11557\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__11580\,
            I => \uu2.un1_w_addr_displaying_inv_4_0\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__11575\,
            I => \uu2.un1_w_addr_displaying_inv_4_0\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__11572\,
            I => \uu2.un1_w_addr_displaying_inv_4_0\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__11569\,
            I => \uu2.un1_w_addr_displaying_inv_4_0\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__11562\,
            I => \uu2.un1_w_addr_displaying_inv_4_0\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__11557\,
            I => \uu2.un1_w_addr_displaying_inv_4_0\
        );

    \I__2274\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11541\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__11541\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_43\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__11538\,
            I => \uu2.segment3_m_1Z0Z_6_cascade_\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__11535\,
            I => \uu2.segment3_m_2_6_cascade_\
        );

    \I__2270\ : InMux
    port map (
            O => \N__11532\,
            I => \N__11529\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__11529\,
            I => \uu2.un1_segment4_4_bmZ0\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__11526\,
            I => \uu2.un1_segment4_4_amZ0_cascade_\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__11523\,
            I => \uu2.N_111_cascade_\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__11520\,
            I => \uu2.un1_segment4_sn_N_36_mux_0_cascade_\
        );

    \I__2265\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11514\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__11514\,
            I => \N__11511\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__11511\,
            I => \uu2.gZ0Z1\
        );

    \I__2262\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11505\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__11505\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_54\
        );

    \I__2260\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11499\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__11499\,
            I => \uu2.un1_segment4_sn_N_58_0\
        );

    \I__2258\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11493\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__11493\,
            I => \uu2.N_2150_0\
        );

    \I__2256\ : InMux
    port map (
            O => \N__11490\,
            I => \N__11487\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__11487\,
            I => \N__11484\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__11484\,
            I => \uu2.un1_segment4_sn_N_38_0_0\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__11481\,
            I => \uu2.g2_1_cascade_\
        );

    \I__2252\ : InMux
    port map (
            O => \N__11478\,
            I => \N__11475\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__11475\,
            I => \N__11472\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__11472\,
            I => \uu2.N_299_0\
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__11469\,
            I => \uu2.g0_i_o4_0_a8_2_2_cascade_\
        );

    \I__2248\ : InMux
    port map (
            O => \N__11466\,
            I => \N__11463\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__11463\,
            I => \uu2.w_addr_displaying_5_rep1_RNIVO2EZ0Z1\
        );

    \I__2246\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11457\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__11457\,
            I => \N__11454\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__11454\,
            I => \uu2.N_315_1_0\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__11451\,
            I => \N__11448\
        );

    \I__2242\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11445\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__11445\,
            I => \uu2.N_94\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__11442\,
            I => \uu2.bitmap_pmux_1_1_3_tz_1_cascade_\
        );

    \I__2239\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11436\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__11436\,
            I => \N__11432\
        );

    \I__2237\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11429\
        );

    \I__2236\ : Span4Mux_h
    port map (
            O => \N__11432\,
            I => \N__11426\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__11429\,
            I => \N__11423\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__11426\,
            I => \uu2.bitmap_pmux_1_1_3_tz\
        );

    \I__2233\ : Odrv12
    port map (
            O => \N__11423\,
            I => \uu2.bitmap_pmux_1_1_3_tz\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__11418\,
            I => \N__11415\
        );

    \I__2231\ : InMux
    port map (
            O => \N__11415\,
            I => \N__11412\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__11412\,
            I => \Lab_UT.didpuu0.didpmtens.N_122\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__11409\,
            I => \N_84_cascade_\
        );

    \I__2228\ : InMux
    port map (
            O => \N__11406\,
            I => \N__11402\
        );

    \I__2227\ : InMux
    port map (
            O => \N__11405\,
            I => \N__11399\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__11402\,
            I => \N_7\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__11399\,
            I => \N_7\
        );

    \I__2224\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11391\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__11391\,
            I => \uu2.un1_segment4_0_bmZ0\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__11388\,
            I => \uu2.un1_segment4_0_amZ0_cascade_\
        );

    \I__2221\ : InMux
    port map (
            O => \N__11385\,
            I => \N__11382\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__11382\,
            I => \N__11379\
        );

    \I__2219\ : Span4Mux_v
    port map (
            O => \N__11379\,
            I => \N__11376\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__11376\,
            I => \uu2.un1_segment4_2_bmZ0\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__11373\,
            I => \uu2.un1_segment4_8_ns_1_cascade_\
        );

    \I__2216\ : InMux
    port map (
            O => \N__11370\,
            I => \N__11367\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__11367\,
            I => \uu2.un1_segment4_2_amZ0\
        );

    \I__2214\ : InMux
    port map (
            O => \N__11364\,
            I => \N__11361\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__11361\,
            I => \uu2.N_286\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__11358\,
            I => \Lab_UT.N_10_cascade_\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__11355\,
            I => \vbuf_tx_data_rdy_cascade_\
        );

    \I__2210\ : CEMux
    port map (
            O => \N__11352\,
            I => \N__11349\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__11349\,
            I => \N__11345\
        );

    \I__2208\ : CEMux
    port map (
            O => \N__11348\,
            I => \N__11342\
        );

    \I__2207\ : Span4Mux_s3_h
    port map (
            O => \N__11345\,
            I => \N__11336\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__11342\,
            I => \N__11336\
        );

    \I__2205\ : CEMux
    port map (
            O => \N__11341\,
            I => \N__11333\
        );

    \I__2204\ : Span4Mux_v
    port map (
            O => \N__11336\,
            I => \N__11328\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__11333\,
            I => \N__11328\
        );

    \I__2202\ : Span4Mux_h
    port map (
            O => \N__11328\,
            I => \N__11325\
        );

    \I__2201\ : Odrv4
    port map (
            O => \N__11325\,
            I => \uu2.vbuf_tx_data_rdy_0\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__11322\,
            I => \N__11319\
        );

    \I__2199\ : InMux
    port map (
            O => \N__11319\,
            I => \N__11316\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__11316\,
            I => \N__11311\
        );

    \I__2197\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11306\
        );

    \I__2196\ : InMux
    port map (
            O => \N__11314\,
            I => \N__11306\
        );

    \I__2195\ : Span4Mux_v
    port map (
            O => \N__11311\,
            I => \N__11299\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__11306\,
            I => \N__11299\
        );

    \I__2193\ : InMux
    port map (
            O => \N__11305\,
            I => \N__11296\
        );

    \I__2192\ : InMux
    port map (
            O => \N__11304\,
            I => \N__11293\
        );

    \I__2191\ : Span4Mux_v
    port map (
            O => \N__11299\,
            I => \N__11290\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__11296\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__11293\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__11290\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__11283\,
            I => \N__11280\
        );

    \I__2186\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11276\
        );

    \I__2185\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11273\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__11276\,
            I => \N__11269\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__11273\,
            I => \N__11266\
        );

    \I__2182\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11263\
        );

    \I__2181\ : Span4Mux_v
    port map (
            O => \N__11269\,
            I => \N__11256\
        );

    \I__2180\ : Span4Mux_v
    port map (
            O => \N__11266\,
            I => \N__11256\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__11263\,
            I => \N__11256\
        );

    \I__2178\ : Span4Mux_h
    port map (
            O => \N__11256\,
            I => \N__11250\
        );

    \I__2177\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11247\
        );

    \I__2176\ : InMux
    port map (
            O => \N__11254\,
            I => \N__11242\
        );

    \I__2175\ : InMux
    port map (
            O => \N__11253\,
            I => \N__11242\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__11250\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__11247\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__11242\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__2171\ : CEMux
    port map (
            O => \N__11235\,
            I => \N__11229\
        );

    \I__2170\ : InMux
    port map (
            O => \N__11234\,
            I => \N__11216\
        );

    \I__2169\ : InMux
    port map (
            O => \N__11233\,
            I => \N__11216\
        );

    \I__2168\ : SRMux
    port map (
            O => \N__11232\,
            I => \N__11213\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__11229\,
            I => \N__11210\
        );

    \I__2166\ : InMux
    port map (
            O => \N__11228\,
            I => \N__11193\
        );

    \I__2165\ : InMux
    port map (
            O => \N__11227\,
            I => \N__11193\
        );

    \I__2164\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11193\
        );

    \I__2163\ : InMux
    port map (
            O => \N__11225\,
            I => \N__11193\
        );

    \I__2162\ : InMux
    port map (
            O => \N__11224\,
            I => \N__11193\
        );

    \I__2161\ : InMux
    port map (
            O => \N__11223\,
            I => \N__11193\
        );

    \I__2160\ : InMux
    port map (
            O => \N__11222\,
            I => \N__11193\
        );

    \I__2159\ : InMux
    port map (
            O => \N__11221\,
            I => \N__11193\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__11216\,
            I => \N__11186\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__11213\,
            I => \N__11183\
        );

    \I__2156\ : Span4Mux_v
    port map (
            O => \N__11210\,
            I => \N__11180\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__11193\,
            I => \N__11177\
        );

    \I__2154\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11170\
        );

    \I__2153\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11170\
        );

    \I__2152\ : InMux
    port map (
            O => \N__11190\,
            I => \N__11170\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__11189\,
            I => \N__11167\
        );

    \I__2150\ : Span4Mux_h
    port map (
            O => \N__11186\,
            I => \N__11159\
        );

    \I__2149\ : Span4Mux_v
    port map (
            O => \N__11183\,
            I => \N__11150\
        );

    \I__2148\ : Span4Mux_s3_h
    port map (
            O => \N__11180\,
            I => \N__11150\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__11177\,
            I => \N__11150\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__11170\,
            I => \N__11150\
        );

    \I__2145\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11147\
        );

    \I__2144\ : InMux
    port map (
            O => \N__11166\,
            I => \N__11142\
        );

    \I__2143\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11142\
        );

    \I__2142\ : InMux
    port map (
            O => \N__11164\,
            I => \N__11139\
        );

    \I__2141\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11136\
        );

    \I__2140\ : InMux
    port map (
            O => \N__11162\,
            I => \N__11133\
        );

    \I__2139\ : Span4Mux_v
    port map (
            O => \N__11159\,
            I => \N__11130\
        );

    \I__2138\ : Span4Mux_v
    port map (
            O => \N__11150\,
            I => \N__11127\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__11147\,
            I => \N__11120\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__11142\,
            I => \N__11120\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__11139\,
            I => \N__11120\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__11136\,
            I => vbuf_tx_data_rdy
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__11133\,
            I => vbuf_tx_data_rdy
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__11130\,
            I => vbuf_tx_data_rdy
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__11127\,
            I => vbuf_tx_data_rdy
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__11120\,
            I => vbuf_tx_data_rdy
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__11109\,
            I => \N__11106\
        );

    \I__2128\ : InMux
    port map (
            O => \N__11106\,
            I => \N__11100\
        );

    \I__2127\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11095\
        );

    \I__2126\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11095\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__11103\,
            I => \N__11092\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__11100\,
            I => \N__11087\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__11095\,
            I => \N__11087\
        );

    \I__2122\ : InMux
    port map (
            O => \N__11092\,
            I => \N__11084\
        );

    \I__2121\ : Span4Mux_v
    port map (
            O => \N__11087\,
            I => \N__11081\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__11084\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__11081\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__2118\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11073\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__11073\,
            I => \N__11065\
        );

    \I__2116\ : InMux
    port map (
            O => \N__11072\,
            I => \N__11058\
        );

    \I__2115\ : InMux
    port map (
            O => \N__11071\,
            I => \N__11058\
        );

    \I__2114\ : InMux
    port map (
            O => \N__11070\,
            I => \N__11058\
        );

    \I__2113\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11053\
        );

    \I__2112\ : InMux
    port map (
            O => \N__11068\,
            I => \N__11053\
        );

    \I__2111\ : Span4Mux_h
    port map (
            O => \N__11065\,
            I => \N__11049\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__11058\,
            I => \N__11046\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__11053\,
            I => \N__11037\
        );

    \I__2108\ : InMux
    port map (
            O => \N__11052\,
            I => \N__11034\
        );

    \I__2107\ : Span4Mux_h
    port map (
            O => \N__11049\,
            I => \N__11031\
        );

    \I__2106\ : Span4Mux_h
    port map (
            O => \N__11046\,
            I => \N__11028\
        );

    \I__2105\ : InMux
    port map (
            O => \N__11045\,
            I => \N__11025\
        );

    \I__2104\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11018\
        );

    \I__2103\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11018\
        );

    \I__2102\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11018\
        );

    \I__2101\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11013\
        );

    \I__2100\ : InMux
    port map (
            O => \N__11040\,
            I => \N__11013\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__11037\,
            I => \N__11008\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__11034\,
            I => \N__11008\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__11031\,
            I => \Lab_UT.secuu0.un4_l_count_0\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__11028\,
            I => \Lab_UT.secuu0.un4_l_count_0\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__11025\,
            I => \Lab_UT.secuu0.un4_l_count_0\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__11018\,
            I => \Lab_UT.secuu0.un4_l_count_0\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__11013\,
            I => \Lab_UT.secuu0.un4_l_count_0\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__11008\,
            I => \Lab_UT.secuu0.un4_l_count_0\
        );

    \I__2091\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10992\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__10992\,
            I => \N__10989\
        );

    \I__2089\ : Span4Mux_h
    port map (
            O => \N__10989\,
            I => \N__10985\
        );

    \I__2088\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10982\
        );

    \I__2087\ : Span4Mux_h
    port map (
            O => \N__10985\,
            I => \N__10977\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__10982\,
            I => \N__10977\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__10977\,
            I => \Lab_UT.secuu0.delay_lineZ0Z_0\
        );

    \I__2084\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10971\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__10971\,
            I => \N__10968\
        );

    \I__2082\ : Span4Mux_s3_h
    port map (
            O => \N__10968\,
            I => \N__10965\
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__10965\,
            I => \Lab_UT.secuu0.delay_lineZ0Z_1\
        );

    \I__2080\ : InMux
    port map (
            O => \N__10962\,
            I => \N__10959\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__10959\,
            I => \resetGen.N_117\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__10956\,
            I => \N__10952\
        );

    \I__2077\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10949\
        );

    \I__2076\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10946\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__10949\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__10946\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__10941\,
            I => \resetGen.N_117_cascade_\
        );

    \I__2072\ : InMux
    port map (
            O => \N__10938\,
            I => \N__10935\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__10935\,
            I => \N__10932\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__10932\,
            I => \N__10928\
        );

    \I__2069\ : IoInMux
    port map (
            O => \N__10931\,
            I => \N__10925\
        );

    \I__2068\ : IoSpan4Mux
    port map (
            O => \N__10928\,
            I => \N__10920\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__10925\,
            I => \N__10920\
        );

    \I__2066\ : IoSpan4Mux
    port map (
            O => \N__10920\,
            I => \N__10917\
        );

    \I__2065\ : Span4Mux_s3_h
    port map (
            O => \N__10917\,
            I => \N__10914\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__10914\,
            I => rst
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__10911\,
            I => \N__10908\
        );

    \I__2062\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10896\
        );

    \I__2061\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10896\
        );

    \I__2060\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10896\
        );

    \I__2059\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10896\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__10896\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__2057\ : InMux
    port map (
            O => \N__10893\,
            I => \N__10884\
        );

    \I__2056\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10884\
        );

    \I__2055\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10884\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__10884\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__2053\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10873\
        );

    \I__2052\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10868\
        );

    \I__2051\ : InMux
    port map (
            O => \N__10879\,
            I => \N__10868\
        );

    \I__2050\ : InMux
    port map (
            O => \N__10878\,
            I => \N__10861\
        );

    \I__2049\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10861\
        );

    \I__2048\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10861\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__10873\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__10868\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__10861\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__10854\,
            I => \resetGen.N_96_cascade_\
        );

    \I__2043\ : InMux
    port map (
            O => \N__10851\,
            I => \N__10839\
        );

    \I__2042\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10839\
        );

    \I__2041\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10839\
        );

    \I__2040\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10839\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__10839\,
            I => \N__10835\
        );

    \I__2038\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10832\
        );

    \I__2037\ : Span4Mux_h
    port map (
            O => \N__10835\,
            I => \N__10829\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__10832\,
            I => \resetGen.N_133\
        );

    \I__2035\ : Odrv4
    port map (
            O => \N__10829\,
            I => \resetGen.N_133\
        );

    \I__2034\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10818\
        );

    \I__2033\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10818\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__10818\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__2031\ : InMux
    port map (
            O => \N__10815\,
            I => \N__10808\
        );

    \I__2030\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10805\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__10813\,
            I => \N__10802\
        );

    \I__2028\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10798\
        );

    \I__2027\ : InMux
    port map (
            O => \N__10811\,
            I => \N__10795\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__10808\,
            I => \N__10790\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__10805\,
            I => \N__10790\
        );

    \I__2024\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10785\
        );

    \I__2023\ : InMux
    port map (
            O => \N__10801\,
            I => \N__10785\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__10798\,
            I => \buart__tx_uart_busy_0\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__10795\,
            I => \buart__tx_uart_busy_0\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__10790\,
            I => \buart__tx_uart_busy_0\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__10785\,
            I => \buart__tx_uart_busy_0\
        );

    \I__2018\ : InMux
    port map (
            O => \N__10776\,
            I => \buart.Z_tx.un1_bitcount_cry_0\
        );

    \I__2017\ : InMux
    port map (
            O => \N__10773\,
            I => \buart.Z_tx.un1_bitcount_cry_1\
        );

    \I__2016\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10767\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__10767\,
            I => \buart.Z_tx.un1_bitcount_axb_3\
        );

    \I__2014\ : InMux
    port map (
            O => \N__10764\,
            I => \buart.Z_tx.un1_bitcount_cry_2\
        );

    \I__2013\ : InMux
    port map (
            O => \N__10761\,
            I => \N__10758\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__10758\,
            I => \buart.Z_tx.bitcount_RNIM5O32Z0Z_2\
        );

    \I__2011\ : InMux
    port map (
            O => \N__10755\,
            I => \N__10752\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__10752\,
            I => \buart.Z_tx.bitcount_RNIL4O32Z0Z_1\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__10749\,
            I => \N__10745\
        );

    \I__2008\ : InMux
    port map (
            O => \N__10748\,
            I => \N__10741\
        );

    \I__2007\ : InMux
    port map (
            O => \N__10745\,
            I => \N__10736\
        );

    \I__2006\ : InMux
    port map (
            O => \N__10744\,
            I => \N__10736\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__10741\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__10736\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__10731\,
            I => \N__10727\
        );

    \I__2002\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10719\
        );

    \I__2001\ : InMux
    port map (
            O => \N__10727\,
            I => \N__10719\
        );

    \I__2000\ : InMux
    port map (
            O => \N__10726\,
            I => \N__10719\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__10719\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__10716\,
            I => \N__10712\
        );

    \I__1997\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10709\
        );

    \I__1996\ : InMux
    port map (
            O => \N__10712\,
            I => \N__10706\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__10709\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__10706\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__10701\,
            I => \N__10697\
        );

    \I__1992\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10692\
        );

    \I__1991\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10689\
        );

    \I__1990\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10684\
        );

    \I__1989\ : InMux
    port map (
            O => \N__10695\,
            I => \N__10684\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__10692\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__10689\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__10684\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__10677\,
            I => \buart__tx_uart_busy_0_cascade_\
        );

    \I__1984\ : InMux
    port map (
            O => \N__10674\,
            I => \N__10663\
        );

    \I__1983\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10656\
        );

    \I__1982\ : InMux
    port map (
            O => \N__10672\,
            I => \N__10656\
        );

    \I__1981\ : InMux
    port map (
            O => \N__10671\,
            I => \N__10656\
        );

    \I__1980\ : InMux
    port map (
            O => \N__10670\,
            I => \N__10651\
        );

    \I__1979\ : InMux
    port map (
            O => \N__10669\,
            I => \N__10651\
        );

    \I__1978\ : InMux
    port map (
            O => \N__10668\,
            I => \N__10644\
        );

    \I__1977\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10644\
        );

    \I__1976\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10644\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__10663\,
            I => \N__10641\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__10656\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__10651\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__10644\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__10641\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1970\ : InMux
    port map (
            O => \N__10632\,
            I => \N__10629\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__10629\,
            I => \buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__10626\,
            I => \N__10623\
        );

    \I__1967\ : InMux
    port map (
            O => \N__10623\,
            I => \N__10620\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__10620\,
            I => \N__10617\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__10617\,
            I => \uu2.un1_segment4_5_bmZ0\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__10614\,
            I => \Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMUZ0Z_0_cascade_\
        );

    \I__1963\ : IoInMux
    port map (
            O => \N__10611\,
            I => \N__10608\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__10608\,
            I => \N__10605\
        );

    \I__1961\ : Span4Mux_s2_h
    port map (
            O => \N__10605\,
            I => \N__10602\
        );

    \I__1960\ : Span4Mux_h
    port map (
            O => \N__10602\,
            I => \N__10599\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__10599\,
            I => led_c_2
        );

    \I__1958\ : InMux
    port map (
            O => \N__10596\,
            I => \N__10593\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__10593\,
            I => \Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJZ0Z_0\
        );

    \I__1956\ : InMux
    port map (
            O => \N__10590\,
            I => \N__10587\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__10587\,
            I => \N__10584\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__10584\,
            I => \uu2.un1_segment4_5_amZ0Z_1\
        );

    \I__1953\ : InMux
    port map (
            O => \N__10581\,
            I => \N__10578\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__10578\,
            I => \uu2.w_addr_displaying_fast_RNIV5694Z0Z_2\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__10575\,
            I => \uu2.N_290_0_i_0_cascade_\
        );

    \I__1950\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10569\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__10569\,
            I => \uu2.w_addr_displaying_RNI362A1Z0Z_3\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__10566\,
            I => \uu2.un1_w_addr_displaying_19_cascade_\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__10563\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_\
        );

    \I__1946\ : InMux
    port map (
            O => \N__10560\,
            I => \N__10557\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__10557\,
            I => \N__10554\
        );

    \I__1944\ : Span4Mux_h
    port map (
            O => \N__10554\,
            I => \N__10551\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__10551\,
            I => \uu2.mem0.N_5_0\
        );

    \I__1942\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10543\
        );

    \I__1941\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10540\
        );

    \I__1940\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10537\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__10543\,
            I => \N__10532\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__10540\,
            I => \N__10532\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__10537\,
            I => \uu2.un1_segment3_s_0\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__10532\,
            I => \uu2.un1_segment3_s_0\
        );

    \I__1935\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10523\
        );

    \I__1934\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10520\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__10523\,
            I => \uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__10520\,
            I => \uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4\
        );

    \I__1931\ : InMux
    port map (
            O => \N__10515\,
            I => \N__10512\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__10512\,
            I => \uu2.mem0.un1_segment3_m2_2\
        );

    \I__1929\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10506\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__10506\,
            I => \uu2.mem0.un1_segment3_m2_0\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__10503\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_42_cascade_\
        );

    \I__1926\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10497\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__10497\,
            I => \N__10494\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__10494\,
            I => \uu2.mem0.un1_segment3_1_0\
        );

    \I__1923\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10488\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__10488\,
            I => \N__10485\
        );

    \I__1921\ : Span4Mux_v
    port map (
            O => \N__10485\,
            I => \N__10482\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__10482\,
            I => \Lab_UT.didpuu0.didpmtens.q_5_0_0_2\
        );

    \I__1919\ : InMux
    port map (
            O => \N__10479\,
            I => \N__10476\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__10476\,
            I => \N__10473\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__10473\,
            I => \uu2.un1_segment4_1_amZ0\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__10470\,
            I => \uu2.un1_segment4_1_bmZ0_cascade_\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__10467\,
            I => \uu2.w_addr_displaying_fast_RNIPN54Z0Z_8_cascade_\
        );

    \I__1914\ : InMux
    port map (
            O => \N__10464\,
            I => \N__10461\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__10461\,
            I => \N__10458\
        );

    \I__1912\ : Odrv4
    port map (
            O => \N__10458\,
            I => \uu2.N_292\
        );

    \I__1911\ : InMux
    port map (
            O => \N__10455\,
            I => \N__10451\
        );

    \I__1910\ : InMux
    port map (
            O => \N__10454\,
            I => \N__10448\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__10451\,
            I => \uu2.N_93\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__10448\,
            I => \uu2.N_93\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__10443\,
            I => \uu2.N_49_cascade_\
        );

    \I__1906\ : InMux
    port map (
            O => \N__10440\,
            I => \N__10437\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__10437\,
            I => \uu2.un1_segment3_m4_s_2\
        );

    \I__1904\ : InMux
    port map (
            O => \N__10434\,
            I => \N__10431\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__10431\,
            I => \uu2.g0_i_o4_0_1\
        );

    \I__1902\ : InMux
    port map (
            O => \N__10428\,
            I => \N__10425\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__10425\,
            I => \uu2.un1_segment3_m4_ns_1\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__10422\,
            I => \uu2.g0_i_o4_3_cascade_\
        );

    \I__1899\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10415\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__10418\,
            I => \N__10410\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__10415\,
            I => \N__10407\
        );

    \I__1896\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10400\
        );

    \I__1895\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10400\
        );

    \I__1894\ : InMux
    port map (
            O => \N__10410\,
            I => \N__10400\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__10407\,
            I => \uu2.un1_segment3_m4\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__10400\,
            I => \uu2.un1_segment3_m4\
        );

    \I__1891\ : InMux
    port map (
            O => \N__10395\,
            I => \N__10392\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__10392\,
            I => \uu2.w_addr_displaying_4_rep1_RNIMMRIAZ0\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__10389\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_53_cascade_\
        );

    \I__1888\ : InMux
    port map (
            O => \N__10386\,
            I => \N__10383\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__10383\,
            I => \uu2.mem0.un1_segment3_1_2\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__10380\,
            I => \Lab_UT_dec3_segmentUQ_1_1_cascade_\
        );

    \I__1885\ : InMux
    port map (
            O => \N__10377\,
            I => \N__10374\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__10374\,
            I => \uu2.Z_decfrac105_7_2\
        );

    \I__1883\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10366\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__10370\,
            I => \N__10361\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__10369\,
            I => \N__10358\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__10366\,
            I => \N__10355\
        );

    \I__1879\ : InMux
    port map (
            O => \N__10365\,
            I => \N__10350\
        );

    \I__1878\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10350\
        );

    \I__1877\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10347\
        );

    \I__1876\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10344\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__10355\,
            I => \N__10339\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__10350\,
            I => \N__10339\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__10347\,
            I => \N__10336\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__10344\,
            I => \N__10333\
        );

    \I__1871\ : Span4Mux_h
    port map (
            O => \N__10339\,
            I => \N__10330\
        );

    \I__1870\ : Span4Mux_v
    port map (
            O => \N__10336\,
            I => \N__10325\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__10333\,
            I => \N__10325\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__10330\,
            I => \Lab_UT.rx_data_0\
        );

    \I__1867\ : Odrv4
    port map (
            O => \N__10325\,
            I => \Lab_UT.rx_data_0\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__10320\,
            I => \N__10317\
        );

    \I__1865\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10313\
        );

    \I__1864\ : InMux
    port map (
            O => \N__10316\,
            I => \N__10309\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__10313\,
            I => \N__10306\
        );

    \I__1862\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10303\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__10309\,
            I => \N__10298\
        );

    \I__1860\ : Span4Mux_v
    port map (
            O => \N__10306\,
            I => \N__10298\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__10303\,
            I => \N__10294\
        );

    \I__1858\ : Span4Mux_h
    port map (
            O => \N__10298\,
            I => \N__10291\
        );

    \I__1857\ : InMux
    port map (
            O => \N__10297\,
            I => \N__10288\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__10294\,
            I => \Lab_UT.rx_dataZ0Z_2\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__10291\,
            I => \Lab_UT.rx_dataZ0Z_2\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__10288\,
            I => \Lab_UT.rx_dataZ0Z_2\
        );

    \I__1853\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10278\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__10278\,
            I => \Lab_UT.dictrluu0.N_103_1\
        );

    \I__1851\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10272\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__10272\,
            I => \N__10269\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__10269\,
            I => \Lab_UT.dicSelectLEDdisp\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__10266\,
            I => \Lab_UT.dicSelectLEDdisp_cascade_\
        );

    \I__1847\ : InMux
    port map (
            O => \N__10263\,
            I => \N__10257\
        );

    \I__1846\ : InMux
    port map (
            O => \N__10262\,
            I => \N__10257\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__10257\,
            I => \N__10254\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__10254\,
            I => \Lab_UT.dictrluu0.N_72\
        );

    \I__1843\ : InMux
    port map (
            O => \N__10251\,
            I => \N__10248\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__10248\,
            I => \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_o2_2\
        );

    \I__1841\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10242\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__10242\,
            I => \N__10239\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__10239\,
            I => \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_3\
        );

    \I__1838\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10233\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__10233\,
            I => \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_4\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__10230\,
            I => \Lab_UT.dictrluu0.dicfsm.N_102_cascade_\
        );

    \I__1835\ : InMux
    port map (
            O => \N__10227\,
            I => \N__10219\
        );

    \I__1834\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10219\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__10225\,
            I => \N__10216\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__10224\,
            I => \N__10213\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__10219\,
            I => \N__10210\
        );

    \I__1830\ : InMux
    port map (
            O => \N__10216\,
            I => \N__10207\
        );

    \I__1829\ : InMux
    port map (
            O => \N__10213\,
            I => \N__10204\
        );

    \I__1828\ : Odrv12
    port map (
            O => \N__10210\,
            I => \Lab_UT_rx_data_7\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__10207\,
            I => \Lab_UT_rx_data_7\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__10204\,
            I => \Lab_UT_rx_data_7\
        );

    \I__1825\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10192\
        );

    \I__1824\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10187\
        );

    \I__1823\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10187\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__10192\,
            I => \N__10184\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__10187\,
            I => \N__10179\
        );

    \I__1820\ : Span4Mux_s3_h
    port map (
            O => \N__10184\,
            I => \N__10176\
        );

    \I__1819\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10171\
        );

    \I__1818\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10171\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__10179\,
            I => \Lab_UT_rx_data_1\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__10176\,
            I => \Lab_UT_rx_data_1\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__10171\,
            I => \Lab_UT_rx_data_1\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__10164\,
            I => \N__10160\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__10163\,
            I => \N__10156\
        );

    \I__1812\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10150\
        );

    \I__1811\ : InMux
    port map (
            O => \N__10159\,
            I => \N__10150\
        );

    \I__1810\ : InMux
    port map (
            O => \N__10156\,
            I => \N__10147\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__10155\,
            I => \N__10144\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__10150\,
            I => \N__10141\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__10147\,
            I => \N__10138\
        );

    \I__1806\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10135\
        );

    \I__1805\ : Odrv12
    port map (
            O => \N__10141\,
            I => \Lab_UT_rx_data_6\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__10138\,
            I => \Lab_UT_rx_data_6\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__10135\,
            I => \Lab_UT_rx_data_6\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__10128\,
            I => \N__10124\
        );

    \I__1801\ : InMux
    port map (
            O => \N__10127\,
            I => \N__10119\
        );

    \I__1800\ : InMux
    port map (
            O => \N__10124\,
            I => \N__10119\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__10119\,
            I => \Lab_UT.rx_data_rdy\
        );

    \I__1798\ : InMux
    port map (
            O => \N__10116\,
            I => \N__10106\
        );

    \I__1797\ : InMux
    port map (
            O => \N__10115\,
            I => \N__10106\
        );

    \I__1796\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10100\
        );

    \I__1795\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10100\
        );

    \I__1794\ : InMux
    port map (
            O => \N__10112\,
            I => \N__10097\
        );

    \I__1793\ : InMux
    port map (
            O => \N__10111\,
            I => \N__10094\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__10106\,
            I => \N__10091\
        );

    \I__1791\ : InMux
    port map (
            O => \N__10105\,
            I => \N__10088\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__10100\,
            I => \N__10085\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__10097\,
            I => \buart__rx_bitcount_0\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__10094\,
            I => \buart__rx_bitcount_0\
        );

    \I__1787\ : Odrv4
    port map (
            O => \N__10091\,
            I => \buart__rx_bitcount_0\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__10088\,
            I => \buart__rx_bitcount_0\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__10085\,
            I => \buart__rx_bitcount_0\
        );

    \I__1784\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10064\
        );

    \I__1783\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10064\
        );

    \I__1782\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10060\
        );

    \I__1781\ : InMux
    port map (
            O => \N__10071\,
            I => \N__10055\
        );

    \I__1780\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10055\
        );

    \I__1779\ : InMux
    port map (
            O => \N__10069\,
            I => \N__10052\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__10064\,
            I => \N__10049\
        );

    \I__1777\ : InMux
    port map (
            O => \N__10063\,
            I => \N__10046\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__10060\,
            I => \N__10043\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__10055\,
            I => \buart__rx_bitcount_2\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__10052\,
            I => \buart__rx_bitcount_2\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__10049\,
            I => \buart__rx_bitcount_2\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__10046\,
            I => \buart__rx_bitcount_2\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__10043\,
            I => \buart__rx_bitcount_2\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__10032\,
            I => \N__10027\
        );

    \I__1769\ : CascadeMux
    port map (
            O => \N__10031\,
            I => \N__10024\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__10030\,
            I => \N__10020\
        );

    \I__1767\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10015\
        );

    \I__1766\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10015\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__10023\,
            I => \N__10010\
        );

    \I__1764\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10006\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__10015\,
            I => \N__10003\
        );

    \I__1762\ : InMux
    port map (
            O => \N__10014\,
            I => \N__10000\
        );

    \I__1761\ : InMux
    port map (
            O => \N__10013\,
            I => \N__9997\
        );

    \I__1760\ : InMux
    port map (
            O => \N__10010\,
            I => \N__9994\
        );

    \I__1759\ : InMux
    port map (
            O => \N__10009\,
            I => \N__9991\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__10006\,
            I => \N__9988\
        );

    \I__1757\ : Span4Mux_h
    port map (
            O => \N__10003\,
            I => \N__9985\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__10000\,
            I => \buart__rx_bitcount_3\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__9997\,
            I => \buart__rx_bitcount_3\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__9994\,
            I => \buart__rx_bitcount_3\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__9991\,
            I => \buart__rx_bitcount_3\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__9988\,
            I => \buart__rx_bitcount_3\
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__9985\,
            I => \buart__rx_bitcount_3\
        );

    \I__1750\ : InMux
    port map (
            O => \N__9972\,
            I => \N__9964\
        );

    \I__1749\ : InMux
    port map (
            O => \N__9971\,
            I => \N__9964\
        );

    \I__1748\ : InMux
    port map (
            O => \N__9970\,
            I => \N__9961\
        );

    \I__1747\ : InMux
    port map (
            O => \N__9969\,
            I => \N__9958\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__9964\,
            I => \N__9955\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__9961\,
            I => \N__9952\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__9958\,
            I => \N_118\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__9955\,
            I => \N_118\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__9952\,
            I => \N_118\
        );

    \I__1741\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9939\
        );

    \I__1740\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9939\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__9939\,
            I => bu_rx_data_rdy
        );

    \I__1738\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9931\
        );

    \I__1737\ : InMux
    port map (
            O => \N__9935\,
            I => \N__9925\
        );

    \I__1736\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9925\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__9931\,
            I => \N__9922\
        );

    \I__1734\ : InMux
    port map (
            O => \N__9930\,
            I => \N__9919\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__9925\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1732\ : Odrv12
    port map (
            O => \N__9922\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__9919\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__1730\ : InMux
    port map (
            O => \N__9912\,
            I => \N__9908\
        );

    \I__1729\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9905\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__9908\,
            I => \buart.Z_rx.N_129\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__9905\,
            I => \buart.Z_rx.N_129\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__9900\,
            I => \bu_rx_data_rdy_cascade_\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__9897\,
            I => \N__9893\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__9896\,
            I => \N__9890\
        );

    \I__1723\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9885\
        );

    \I__1722\ : InMux
    port map (
            O => \N__9890\,
            I => \N__9880\
        );

    \I__1721\ : InMux
    port map (
            O => \N__9889\,
            I => \N__9880\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__9888\,
            I => \N__9876\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__9885\,
            I => \N__9865\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__9880\,
            I => \N__9865\
        );

    \I__1717\ : InMux
    port map (
            O => \N__9879\,
            I => \N__9862\
        );

    \I__1716\ : InMux
    port map (
            O => \N__9876\,
            I => \N__9853\
        );

    \I__1715\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9853\
        );

    \I__1714\ : InMux
    port map (
            O => \N__9874\,
            I => \N__9853\
        );

    \I__1713\ : InMux
    port map (
            O => \N__9873\,
            I => \N__9853\
        );

    \I__1712\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9846\
        );

    \I__1711\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9846\
        );

    \I__1710\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9846\
        );

    \I__1709\ : Span4Mux_s3_v
    port map (
            O => \N__9865\,
            I => \N__9842\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__9862\,
            I => \N__9835\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__9853\,
            I => \N__9835\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__9846\,
            I => \N__9835\
        );

    \I__1705\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9832\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__9842\,
            I => \buart.Z_rx.startbit\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__9835\,
            I => \buart.Z_rx.startbit\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__9832\,
            I => \buart.Z_rx.startbit\
        );

    \I__1701\ : CEMux
    port map (
            O => \N__9825\,
            I => \N__9821\
        );

    \I__1700\ : CEMux
    port map (
            O => \N__9824\,
            I => \N__9818\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__9821\,
            I => \N__9815\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__9818\,
            I => \N__9812\
        );

    \I__1697\ : Span4Mux_s3_v
    port map (
            O => \N__9815\,
            I => \N__9807\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__9812\,
            I => \N__9807\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__9807\,
            I => \buart.Z_rx.bitcount_e_0_RNII0231Z0Z_0\
        );

    \I__1694\ : CascadeMux
    port map (
            O => \N__9804\,
            I => \Lab_UT_dec3_segmentUQ_0_6_cascade_\
        );

    \I__1693\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9798\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__9798\,
            I => \N_71\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__9795\,
            I => \N_71_cascade_\
        );

    \I__1690\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9785\
        );

    \I__1689\ : InMux
    port map (
            O => \N__9791\,
            I => \N__9785\
        );

    \I__1688\ : InMux
    port map (
            O => \N__9790\,
            I => \N__9782\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__9785\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__9782\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__1685\ : InMux
    port map (
            O => \N__9777\,
            I => \N__9773\
        );

    \I__1684\ : InMux
    port map (
            O => \N__9776\,
            I => \N__9770\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__9773\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__9770\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__9765\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__9762\,
            I => \N__9756\
        );

    \I__1679\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9749\
        );

    \I__1678\ : InMux
    port map (
            O => \N__9760\,
            I => \N__9749\
        );

    \I__1677\ : InMux
    port map (
            O => \N__9759\,
            I => \N__9749\
        );

    \I__1676\ : InMux
    port map (
            O => \N__9756\,
            I => \N__9746\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__9749\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__9746\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__1673\ : InMux
    port map (
            O => \N__9741\,
            I => \N__9738\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__9738\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__9735\,
            I => \buart.Z_rx.ser_clk_cascade_\
        );

    \I__1670\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9727\
        );

    \I__1669\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9722\
        );

    \I__1668\ : InMux
    port map (
            O => \N__9730\,
            I => \N__9722\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__9727\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__9722\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__1665\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9714\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__9714\,
            I => \N__9710\
        );

    \I__1663\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9706\
        );

    \I__1662\ : Span4Mux_h
    port map (
            O => \N__9710\,
            I => \N__9703\
        );

    \I__1661\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9700\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__9706\,
            I => \N__9697\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__9703\,
            I => bu_rx_data_7
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__9700\,
            I => bu_rx_data_7
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__9697\,
            I => bu_rx_data_7
        );

    \I__1656\ : InMux
    port map (
            O => \N__9690\,
            I => \N__9687\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__9687\,
            I => \N__9683\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__9686\,
            I => \N__9679\
        );

    \I__1653\ : Span4Mux_h
    port map (
            O => \N__9683\,
            I => \N__9676\
        );

    \I__1652\ : InMux
    port map (
            O => \N__9682\,
            I => \N__9671\
        );

    \I__1651\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9671\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__9676\,
            I => bu_rx_data_6
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__9671\,
            I => bu_rx_data_6
        );

    \I__1648\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9663\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__9663\,
            I => \N__9660\
        );

    \I__1646\ : Span12Mux_s5_h
    port map (
            O => \N__9660\,
            I => \N__9655\
        );

    \I__1645\ : InMux
    port map (
            O => \N__9659\,
            I => \N__9652\
        );

    \I__1644\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9649\
        );

    \I__1643\ : Odrv12
    port map (
            O => \N__9655\,
            I => bu_rx_data_2
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__9652\,
            I => bu_rx_data_2
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__9649\,
            I => bu_rx_data_2
        );

    \I__1640\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9639\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__9639\,
            I => \N__9636\
        );

    \I__1638\ : Span4Mux_h
    port map (
            O => \N__9636\,
            I => \N__9631\
        );

    \I__1637\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9628\
        );

    \I__1636\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9625\
        );

    \I__1635\ : Odrv4
    port map (
            O => \N__9631\,
            I => bu_rx_data_4
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__9628\,
            I => bu_rx_data_4
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__9625\,
            I => bu_rx_data_4
        );

    \I__1632\ : InMux
    port map (
            O => \N__9618\,
            I => \N__9615\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__9615\,
            I => \N__9611\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__9614\,
            I => \N__9607\
        );

    \I__1629\ : Span4Mux_v
    port map (
            O => \N__9611\,
            I => \N__9604\
        );

    \I__1628\ : InMux
    port map (
            O => \N__9610\,
            I => \N__9601\
        );

    \I__1627\ : InMux
    port map (
            O => \N__9607\,
            I => \N__9598\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__9604\,
            I => bu_rx_data_3
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__9601\,
            I => bu_rx_data_3
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__9598\,
            I => bu_rx_data_3
        );

    \I__1623\ : InMux
    port map (
            O => \N__9591\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__1622\ : InMux
    port map (
            O => \N__9588\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__1621\ : InMux
    port map (
            O => \N__9585\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__1620\ : InMux
    port map (
            O => \N__9582\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__9579\,
            I => \N__9576\
        );

    \I__1618\ : InMux
    port map (
            O => \N__9576\,
            I => \N__9573\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__9573\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__1616\ : CEMux
    port map (
            O => \N__9570\,
            I => \N__9567\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__9567\,
            I => \N__9564\
        );

    \I__1614\ : Span4Mux_v
    port map (
            O => \N__9564\,
            I => \N__9561\
        );

    \I__1613\ : Span4Mux_s0_v
    port map (
            O => \N__9561\,
            I => \N__9557\
        );

    \I__1612\ : CEMux
    port map (
            O => \N__9560\,
            I => \N__9554\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__9557\,
            I => \N__9549\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__9554\,
            I => \N__9549\
        );

    \I__1609\ : Span4Mux_v
    port map (
            O => \N__9549\,
            I => \N__9546\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__9546\,
            I => \N__9543\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__9543\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1606\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9536\
        );

    \I__1605\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9533\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__9536\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__9533\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__9528\,
            I => \N__9523\
        );

    \I__1601\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9520\
        );

    \I__1600\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9515\
        );

    \I__1599\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9515\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__9520\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__9515\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1596\ : InMux
    port map (
            O => \N__9510\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__1595\ : InMux
    port map (
            O => \N__9507\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__1594\ : InMux
    port map (
            O => \N__9504\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__9501\,
            I => \N__9498\
        );

    \I__1592\ : InMux
    port map (
            O => \N__9498\,
            I => \N__9492\
        );

    \I__1591\ : InMux
    port map (
            O => \N__9497\,
            I => \N__9492\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__9492\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__9489\,
            I => \N__9486\
        );

    \I__1588\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9480\
        );

    \I__1587\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9480\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__9480\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__9477\,
            I => \N__9473\
        );

    \I__1584\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9470\
        );

    \I__1583\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9467\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__9470\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__9467\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__9462\,
            I => \N__9459\
        );

    \I__1579\ : InMux
    port map (
            O => \N__9459\,
            I => \N__9453\
        );

    \I__1578\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9453\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__9453\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__9450\,
            I => \N__9446\
        );

    \I__1575\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9441\
        );

    \I__1574\ : InMux
    port map (
            O => \N__9446\,
            I => \N__9441\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__9441\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__1572\ : InMux
    port map (
            O => \N__9438\,
            I => \N__9435\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__9435\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__1570\ : InMux
    port map (
            O => \N__9432\,
            I => \N__9424\
        );

    \I__1569\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9424\
        );

    \I__1568\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9421\
        );

    \I__1567\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9418\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__9424\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__9421\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__9418\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__9411\,
            I => \N__9407\
        );

    \I__1562\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9403\
        );

    \I__1561\ : InMux
    port map (
            O => \N__9407\,
            I => \N__9400\
        );

    \I__1560\ : InMux
    port map (
            O => \N__9406\,
            I => \N__9397\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__9403\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__9400\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__9397\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__1556\ : InMux
    port map (
            O => \N__9390\,
            I => \N__9387\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__9387\,
            I => vbuf_tx_data_7
        );

    \I__1554\ : InMux
    port map (
            O => \N__9384\,
            I => \N__9381\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__9381\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__1552\ : CascadeMux
    port map (
            O => \N__9378\,
            I => \N__9375\
        );

    \I__1551\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9372\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__9372\,
            I => \N__9367\
        );

    \I__1549\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9362\
        );

    \I__1548\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9359\
        );

    \I__1547\ : Span4Mux_h
    port map (
            O => \N__9367\,
            I => \N__9356\
        );

    \I__1546\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9351\
        );

    \I__1545\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9351\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__9362\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__9359\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__9356\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__9351\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__9342\,
            I => \N__9339\
        );

    \I__1539\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9336\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__9336\,
            I => \N__9333\
        );

    \I__1537\ : Span4Mux_h
    port map (
            O => \N__9333\,
            I => \N__9330\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__9330\,
            I => \uu2.mem0.w_addr_4\
        );

    \I__1535\ : InMux
    port map (
            O => \N__9327\,
            I => \N__9324\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__9324\,
            I => \N__9319\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__9323\,
            I => \N__9315\
        );

    \I__1532\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9312\
        );

    \I__1531\ : Span4Mux_h
    port map (
            O => \N__9319\,
            I => \N__9309\
        );

    \I__1530\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9304\
        );

    \I__1529\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9304\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__9312\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__9309\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__9304\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__9297\,
            I => \N__9294\
        );

    \I__1524\ : InMux
    port map (
            O => \N__9294\,
            I => \N__9291\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__9291\,
            I => \N__9288\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__9288\,
            I => \N__9285\
        );

    \I__1521\ : Span4Mux_s2_h
    port map (
            O => \N__9285\,
            I => \N__9282\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__9282\,
            I => \uu2.mem0.w_addr_5\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__9279\,
            I => \N__9276\
        );

    \I__1518\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9273\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__9273\,
            I => \N__9270\
        );

    \I__1516\ : Odrv4
    port map (
            O => \N__9270\,
            I => \uu2.Z_decfrac106_2\
        );

    \I__1515\ : InMux
    port map (
            O => \N__9267\,
            I => \N__9264\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__9264\,
            I => \N__9261\
        );

    \I__1513\ : Span4Mux_h
    port map (
            O => \N__9261\,
            I => \N__9258\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__9258\,
            I => \uu2.mem0.N_2160_1\
        );

    \I__1511\ : InMux
    port map (
            O => \N__9255\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__1510\ : InMux
    port map (
            O => \N__9252\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__1509\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9246\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__9246\,
            I => \uu2.mem0.un1_segment3_0\
        );

    \I__1507\ : InMux
    port map (
            O => \N__9243\,
            I => \N__9240\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__9240\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_34\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__9237\,
            I => \N__9232\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__9236\,
            I => \N__9229\
        );

    \I__1503\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9221\
        );

    \I__1502\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9221\
        );

    \I__1501\ : InMux
    port map (
            O => \N__9229\,
            I => \N__9221\
        );

    \I__1500\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9218\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__9221\,
            I => \N__9212\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__9218\,
            I => \N__9212\
        );

    \I__1497\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9209\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__9212\,
            I => \uu2.Z_decfrac106\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__9209\,
            I => \uu2.Z_decfrac106\
        );

    \I__1494\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9201\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__9201\,
            I => \uu2.mem0.un1_segment3_m2_1\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__9198\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_47_cascade_\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__9195\,
            I => \N__9192\
        );

    \I__1490\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9189\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__9189\,
            I => \uu2.mem0.un1_segment3_1_1\
        );

    \I__1488\ : InMux
    port map (
            O => \N__9186\,
            I => \N__9183\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__9183\,
            I => \uu2.mem0.N_2160_0\
        );

    \I__1486\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9177\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__9177\,
            I => \N__9174\
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__9174\,
            I => \N_52\
        );

    \I__1483\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9168\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__9168\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_48\
        );

    \I__1481\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9162\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__9162\,
            I => vbuf_tx_data_6
        );

    \I__1479\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9156\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__9156\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__1477\ : InMux
    port map (
            O => \N__9153\,
            I => \N__9150\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__9150\,
            I => \N__9147\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__9147\,
            I => \N_52_0\
        );

    \I__1474\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9141\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__9141\,
            I => \L3_segment2_0_0\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__9138\,
            I => \uu2.mem0.N_2159_0_cascade_\
        );

    \I__1471\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9132\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__9132\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_20\
        );

    \I__1469\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9126\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__9126\,
            I => \N__9123\
        );

    \I__1467\ : Odrv12
    port map (
            O => \N__9123\,
            I => \L3_segment2_0\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__9120\,
            I => \uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4_cascade_\
        );

    \I__1465\ : InMux
    port map (
            O => \N__9117\,
            I => \N__9114\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__9114\,
            I => \uu2.mem0.g2_0\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__9111\,
            I => \uu2.mem0.N_5_cascade_\
        );

    \I__1462\ : InMux
    port map (
            O => \N__9108\,
            I => \N__9105\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__9105\,
            I => \uu2.mem0.bitmap_pmux_1_1_0_0\
        );

    \I__1460\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9099\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__9099\,
            I => \uu2.mem0.N_14\
        );

    \I__1458\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9093\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__9093\,
            I => \uu2.mem0.N_18\
        );

    \I__1456\ : CEMux
    port map (
            O => \N__9090\,
            I => \N__9087\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__9087\,
            I => \N__9084\
        );

    \I__1454\ : Span4Mux_s1_h
    port map (
            O => \N__9084\,
            I => \N__9079\
        );

    \I__1453\ : CEMux
    port map (
            O => \N__9083\,
            I => \N__9076\
        );

    \I__1452\ : CEMux
    port map (
            O => \N__9082\,
            I => \N__9073\
        );

    \I__1451\ : Span4Mux_v
    port map (
            O => \N__9079\,
            I => \N__9070\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__9076\,
            I => \N__9067\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__9073\,
            I => \N__9064\
        );

    \I__1448\ : Span4Mux_h
    port map (
            O => \N__9070\,
            I => \N__9061\
        );

    \I__1447\ : Span4Mux_s2_h
    port map (
            O => \N__9067\,
            I => \N__9058\
        );

    \I__1446\ : Span4Mux_h
    port map (
            O => \N__9064\,
            I => \N__9055\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__9061\,
            I => \Lab_UT.Lab3U00.bu_rx_data_rdy_0\
        );

    \I__1444\ : Odrv4
    port map (
            O => \N__9058\,
            I => \Lab_UT.Lab3U00.bu_rx_data_rdy_0\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__9055\,
            I => \Lab_UT.Lab3U00.bu_rx_data_rdy_0\
        );

    \I__1442\ : InMux
    port map (
            O => \N__9048\,
            I => \N__9043\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__9047\,
            I => \N__9040\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__9046\,
            I => \N__9037\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__9043\,
            I => \N__9032\
        );

    \I__1438\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9029\
        );

    \I__1437\ : InMux
    port map (
            O => \N__9037\,
            I => \N__9026\
        );

    \I__1436\ : InMux
    port map (
            O => \N__9036\,
            I => \N__9021\
        );

    \I__1435\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9021\
        );

    \I__1434\ : Span4Mux_h
    port map (
            O => \N__9032\,
            I => \N__9018\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__9029\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__9026\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__9021\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__9018\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__9009\,
            I => \N__9006\
        );

    \I__1428\ : InMux
    port map (
            O => \N__9006\,
            I => \N__9003\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__9003\,
            I => \N__9000\
        );

    \I__1426\ : Span4Mux_v
    port map (
            O => \N__9000\,
            I => \N__8997\
        );

    \I__1425\ : Odrv4
    port map (
            O => \N__8997\,
            I => \uu2.mem0.w_addr_2\
        );

    \I__1424\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8991\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__8991\,
            I => \N__8984\
        );

    \I__1422\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8979\
        );

    \I__1421\ : InMux
    port map (
            O => \N__8989\,
            I => \N__8979\
        );

    \I__1420\ : InMux
    port map (
            O => \N__8988\,
            I => \N__8974\
        );

    \I__1419\ : InMux
    port map (
            O => \N__8987\,
            I => \N__8974\
        );

    \I__1418\ : Span4Mux_h
    port map (
            O => \N__8984\,
            I => \N__8971\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__8979\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__8974\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__8971\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__8964\,
            I => \N__8961\
        );

    \I__1413\ : InMux
    port map (
            O => \N__8961\,
            I => \N__8958\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__8958\,
            I => \N__8955\
        );

    \I__1411\ : Span4Mux_h
    port map (
            O => \N__8955\,
            I => \N__8952\
        );

    \I__1410\ : Odrv4
    port map (
            O => \N__8952\,
            I => \uu2.mem0.w_addr_3\
        );

    \I__1409\ : InMux
    port map (
            O => \N__8949\,
            I => \N__8946\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__8946\,
            I => \uu2.mem0.G_14_0_0\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__8943\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_32_cascade_\
        );

    \I__1406\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8937\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__8937\,
            I => \uu2.mem0.G_14_0_1\
        );

    \I__1404\ : CascadeMux
    port map (
            O => \N__8934\,
            I => \uu2.N_329_0_cascade_\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__8931\,
            I => \N__8928\
        );

    \I__1402\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8923\
        );

    \I__1401\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8920\
        );

    \I__1400\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8914\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__8923\,
            I => \N__8911\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__8920\,
            I => \N__8908\
        );

    \I__1397\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8903\
        );

    \I__1396\ : InMux
    port map (
            O => \N__8918\,
            I => \N__8903\
        );

    \I__1395\ : InMux
    port map (
            O => \N__8917\,
            I => \N__8900\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__8914\,
            I => \N__8897\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__8911\,
            I => \uu2.Z_decfrac105_7\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__8908\,
            I => \uu2.Z_decfrac105_7\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__8903\,
            I => \uu2.Z_decfrac105_7\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__8900\,
            I => \uu2.Z_decfrac105_7\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__8897\,
            I => \uu2.Z_decfrac105_7\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__8886\,
            I => \N__8882\
        );

    \I__1387\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8876\
        );

    \I__1386\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8867\
        );

    \I__1385\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8867\
        );

    \I__1384\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8867\
        );

    \I__1383\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8867\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__8876\,
            I => \N__8862\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__8867\,
            I => \N__8862\
        );

    \I__1380\ : Odrv12
    port map (
            O => \N__8862\,
            I => \buart.Z_rx.N_39\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__8859\,
            I => \N__8854\
        );

    \I__1378\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8849\
        );

    \I__1377\ : InMux
    port map (
            O => \N__8857\,
            I => \N__8849\
        );

    \I__1376\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8846\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__8849\,
            I => \N__8843\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__8846\,
            I => \N__8838\
        );

    \I__1373\ : Span4Mux_v
    port map (
            O => \N__8843\,
            I => \N__8835\
        );

    \I__1372\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8832\
        );

    \I__1371\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8829\
        );

    \I__1370\ : Odrv12
    port map (
            O => \N__8838\,
            I => \Lab_UT_rx_data_4\
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__8835\,
            I => \Lab_UT_rx_data_4\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__8832\,
            I => \Lab_UT_rx_data_4\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__8829\,
            I => \Lab_UT_rx_data_4\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__8820\,
            I => \N__8817\
        );

    \I__1365\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8812\
        );

    \I__1364\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8809\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__8815\,
            I => \N__8805\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__8812\,
            I => \N__8800\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__8809\,
            I => \N__8800\
        );

    \I__1360\ : InMux
    port map (
            O => \N__8808\,
            I => \N__8795\
        );

    \I__1359\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8795\
        );

    \I__1358\ : Span4Mux_h
    port map (
            O => \N__8800\,
            I => \N__8792\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__8795\,
            I => \N__8789\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__8792\,
            I => \Lab_UT_rx_data_3\
        );

    \I__1355\ : Odrv12
    port map (
            O => \N__8789\,
            I => \Lab_UT_rx_data_3\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__8784\,
            I => \Lab_UT.dictrluu0.N_103_1_cascade_\
        );

    \I__1353\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8778\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__8778\,
            I => \N__8775\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__8775\,
            I => \N__8769\
        );

    \I__1350\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8766\
        );

    \I__1349\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8761\
        );

    \I__1348\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8761\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__8769\,
            I => \Lab_UT_rx_data_5\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__8766\,
            I => \Lab_UT_rx_data_5\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__8761\,
            I => \Lab_UT_rx_data_5\
        );

    \I__1344\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8751\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__8751\,
            I => \N__8748\
        );

    \I__1342\ : Odrv12
    port map (
            O => \N__8748\,
            I => \uu2.un1_w_user_lf_3Z0Z_1\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__8745\,
            I => \N__8738\
        );

    \I__1340\ : InMux
    port map (
            O => \N__8744\,
            I => \N__8732\
        );

    \I__1339\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8732\
        );

    \I__1338\ : InMux
    port map (
            O => \N__8742\,
            I => \N__8718\
        );

    \I__1337\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8715\
        );

    \I__1336\ : InMux
    port map (
            O => \N__8738\,
            I => \N__8710\
        );

    \I__1335\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8710\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__8732\,
            I => \N__8707\
        );

    \I__1333\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8700\
        );

    \I__1332\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8700\
        );

    \I__1331\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8700\
        );

    \I__1330\ : InMux
    port map (
            O => \N__8728\,
            I => \N__8693\
        );

    \I__1329\ : InMux
    port map (
            O => \N__8727\,
            I => \N__8693\
        );

    \I__1328\ : InMux
    port map (
            O => \N__8726\,
            I => \N__8693\
        );

    \I__1327\ : InMux
    port map (
            O => \N__8725\,
            I => \N__8682\
        );

    \I__1326\ : InMux
    port map (
            O => \N__8724\,
            I => \N__8682\
        );

    \I__1325\ : InMux
    port map (
            O => \N__8723\,
            I => \N__8682\
        );

    \I__1324\ : InMux
    port map (
            O => \N__8722\,
            I => \N__8682\
        );

    \I__1323\ : InMux
    port map (
            O => \N__8721\,
            I => \N__8682\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__8718\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__8715\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__8710\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__1319\ : Odrv12
    port map (
            O => \N__8707\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__8700\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__8693\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__8682\,
            I => \Lab_UT_dspStr_cnt_1\
        );

    \I__1315\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8661\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__8666\,
            I => \N__8646\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__8665\,
            I => \N__8643\
        );

    \I__1312\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8639\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__8661\,
            I => \N__8636\
        );

    \I__1310\ : InMux
    port map (
            O => \N__8660\,
            I => \N__8633\
        );

    \I__1309\ : InMux
    port map (
            O => \N__8659\,
            I => \N__8628\
        );

    \I__1308\ : InMux
    port map (
            O => \N__8658\,
            I => \N__8628\
        );

    \I__1307\ : InMux
    port map (
            O => \N__8657\,
            I => \N__8625\
        );

    \I__1306\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8620\
        );

    \I__1305\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8620\
        );

    \I__1304\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8613\
        );

    \I__1303\ : InMux
    port map (
            O => \N__8653\,
            I => \N__8613\
        );

    \I__1302\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8613\
        );

    \I__1301\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8606\
        );

    \I__1300\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8606\
        );

    \I__1299\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8606\
        );

    \I__1298\ : InMux
    port map (
            O => \N__8646\,
            I => \N__8599\
        );

    \I__1297\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8599\
        );

    \I__1296\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8599\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__8639\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__1294\ : Odrv12
    port map (
            O => \N__8636\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__8633\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__8628\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__8625\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__8620\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__8613\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__8606\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__8599\,
            I => \Lab_UT_dspStr_cnt_3\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__8580\,
            I => \uu2.mem0.N_26_1_cascade_\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__8577\,
            I => \N__8571\
        );

    \I__1284\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8555\
        );

    \I__1283\ : InMux
    port map (
            O => \N__8575\,
            I => \N__8555\
        );

    \I__1282\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8552\
        );

    \I__1281\ : InMux
    port map (
            O => \N__8571\,
            I => \N__8549\
        );

    \I__1280\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8546\
        );

    \I__1279\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8543\
        );

    \I__1278\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8536\
        );

    \I__1277\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8536\
        );

    \I__1276\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8536\
        );

    \I__1275\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8529\
        );

    \I__1274\ : InMux
    port map (
            O => \N__8564\,
            I => \N__8529\
        );

    \I__1273\ : InMux
    port map (
            O => \N__8563\,
            I => \N__8529\
        );

    \I__1272\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8522\
        );

    \I__1271\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8522\
        );

    \I__1270\ : InMux
    port map (
            O => \N__8560\,
            I => \N__8522\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__8555\,
            I => \N__8519\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__8552\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__8549\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__8546\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__8543\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__8536\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__8529\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__8522\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__1261\ : Odrv12
    port map (
            O => \N__8519\,
            I => \Lab_UT_dspStr_cnt_2\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__8502\,
            I => \resetGen.reset_count_2_i_0_a3_5Z0Z_4_cascade_\
        );

    \I__1259\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8496\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__1257\ : Span4Mux_v
    port map (
            O => \N__8493\,
            I => \N__8488\
        );

    \I__1256\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8483\
        );

    \I__1255\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8483\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__8488\,
            I => bu_rx_data_5
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__8483\,
            I => bu_rx_data_5
        );

    \I__1252\ : InMux
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__8475\,
            I => \resetGen.reset_count_2_i_0_a3_6Z0Z_4\
        );

    \I__1250\ : InMux
    port map (
            O => \N__8472\,
            I => \N__8469\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__8469\,
            I => \resetGen.reset_count_2_i_0_a3_4Z0Z_4\
        );

    \I__1248\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8462\
        );

    \I__1247\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8459\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__8462\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__8459\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__8454\,
            I => \buart.Z_rx.N_129_cascade_\
        );

    \I__1243\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8445\
        );

    \I__1242\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8445\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__8445\,
            I => \N__8442\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__8442\,
            I => \N__8439\
        );

    \I__1239\ : Span4Mux_h
    port map (
            O => \N__8439\,
            I => \N__8436\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__8436\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1237\ : InMux
    port map (
            O => \N__8433\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__8430\,
            I => \buart.Z_rx.N_144_cascade_\
        );

    \I__1235\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8422\
        );

    \I__1234\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8417\
        );

    \I__1233\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8417\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__8422\,
            I => \buart__rx_bitcount_4\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__8417\,
            I => \buart__rx_bitcount_4\
        );

    \I__1230\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8409\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__8409\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__1228\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8400\
        );

    \I__1227\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8397\
        );

    \I__1226\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8392\
        );

    \I__1225\ : InMux
    port map (
            O => \N__8403\,
            I => \N__8392\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__8400\,
            I => \buart__rx_bitcount_1\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__8397\,
            I => \buart__rx_bitcount_1\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__8392\,
            I => \buart__rx_bitcount_1\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__8385\,
            I => \N__8382\
        );

    \I__1220\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8379\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__8379\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__1218\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8373\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__8373\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__1216\ : IoInMux
    port map (
            O => \N__8370\,
            I => \N__8366\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__8369\,
            I => \N__8363\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__8366\,
            I => \N__8360\
        );

    \I__1213\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8357\
        );

    \I__1212\ : Span4Mux_s1_v
    port map (
            O => \N__8360\,
            I => \N__8354\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__8357\,
            I => \N__8351\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__8354\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1209\ : Odrv12
    port map (
            O => \N__8351\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1208\ : InMux
    port map (
            O => \N__8346\,
            I => \N__8343\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__8343\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__1206\ : InMux
    port map (
            O => \N__8340\,
            I => \N__8337\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__8337\,
            I => \N__8334\
        );

    \I__1204\ : Span4Mux_v
    port map (
            O => \N__8334\,
            I => \N__8331\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__8331\,
            I => vbuf_tx_data_3
        );

    \I__1202\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8325\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__8325\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__1200\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8319\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__8319\,
            I => vbuf_tx_data_4
        );

    \I__1198\ : InMux
    port map (
            O => \N__8316\,
            I => \N__8313\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__8313\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__1196\ : InMux
    port map (
            O => \N__8310\,
            I => \N__8307\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__8307\,
            I => vbuf_tx_data_5
        );

    \I__1194\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8301\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__8301\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__1192\ : InMux
    port map (
            O => \N__8298\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__1191\ : InMux
    port map (
            O => \N__8295\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__1190\ : InMux
    port map (
            O => \N__8292\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__1189\ : InMux
    port map (
            O => \N__8289\,
            I => \N__8286\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__8286\,
            I => \N__8283\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__8283\,
            I => \uu2.r_data_wire_4\
        );

    \I__1186\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8277\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__8277\,
            I => \N__8274\
        );

    \I__1184\ : Odrv4
    port map (
            O => \N__8274\,
            I => \uu2.r_data_wire_5\
        );

    \I__1183\ : InMux
    port map (
            O => \N__8271\,
            I => \N__8268\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__8268\,
            I => \N__8265\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__8265\,
            I => \uu2.r_data_wire_6\
        );

    \I__1180\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8259\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__8259\,
            I => \N__8256\
        );

    \I__1178\ : Odrv4
    port map (
            O => \N__8256\,
            I => \uu2.r_data_wire_7\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__8253\,
            I => \N__8250\
        );

    \I__1176\ : InMux
    port map (
            O => \N__8250\,
            I => \N__8247\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__8247\,
            I => vbuf_tx_data_0
        );

    \I__1174\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8241\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__8241\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__1172\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8235\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__8235\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__1170\ : IoInMux
    port map (
            O => \N__8232\,
            I => \N__8229\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__8229\,
            I => \N__8226\
        );

    \I__1168\ : Span4Mux_s3_h
    port map (
            O => \N__8226\,
            I => \N__8223\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__8223\,
            I => o_serial_data_c
        );

    \I__1166\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8217\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__8217\,
            I => vbuf_tx_data_1
        );

    \I__1164\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8211\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__8211\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__1162\ : InMux
    port map (
            O => \N__8208\,
            I => \N__8205\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__8205\,
            I => vbuf_tx_data_2
        );

    \I__1160\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8199\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__8199\,
            I => \uu2.bitmap_pmux_1_1_a8_1_2_0\
        );

    \I__1158\ : InMux
    port map (
            O => \N__8196\,
            I => \N__8193\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__8193\,
            I => \uu2.N_326_0\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__8190\,
            I => \uu2.bitmap_pmux_1_1_a8_1_1_cascade_\
        );

    \I__1155\ : InMux
    port map (
            O => \N__8187\,
            I => \N__8184\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__8184\,
            I => \uu2.bitmap_pmux_1_1_a8_0_1\
        );

    \I__1153\ : InMux
    port map (
            O => \N__8181\,
            I => \N__8178\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__8178\,
            I => \uu2.bitmap_pmux_1_1_1_tz\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__8175\,
            I => \uu2.bitmap_pmux_1_1_1_tz_cascade_\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__8172\,
            I => \N__8169\
        );

    \I__1149\ : InMux
    port map (
            O => \N__8169\,
            I => \N__8166\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__8166\,
            I => \N__8163\
        );

    \I__1147\ : Span4Mux_v
    port map (
            O => \N__8163\,
            I => \N__8159\
        );

    \I__1146\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8156\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__8159\,
            I => \L3_tx_data_3\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__8156\,
            I => \L3_tx_data_3\
        );

    \I__1143\ : InMux
    port map (
            O => \N__8151\,
            I => \N__8148\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__8148\,
            I => \N__8145\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__8145\,
            I => \uu2.mem0.w_data_1_0_0_3\
        );

    \I__1140\ : IoInMux
    port map (
            O => \N__8142\,
            I => \N__8138\
        );

    \I__1139\ : InMux
    port map (
            O => \N__8141\,
            I => \N__8135\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__8138\,
            I => \N__8132\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__8135\,
            I => \N__8129\
        );

    \I__1136\ : Span12Mux_s5_v
    port map (
            O => \N__8132\,
            I => \N__8124\
        );

    \I__1135\ : Span12Mux_s5_h
    port map (
            O => \N__8129\,
            I => \N__8124\
        );

    \I__1134\ : Odrv12
    port map (
            O => \N__8124\,
            I => \latticehx1k_pll_inst_PLLOUTCORE_i\
        );

    \I__1133\ : CEMux
    port map (
            O => \N__8121\,
            I => \N__8117\
        );

    \I__1132\ : SRMux
    port map (
            O => \N__8120\,
            I => \N__8114\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__8117\,
            I => \N__8111\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__8114\,
            I => \N__8108\
        );

    \I__1129\ : Span4Mux_v
    port map (
            O => \N__8111\,
            I => \N__8105\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__8108\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__8105\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1126\ : InMux
    port map (
            O => \N__8100\,
            I => \N__8097\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__8097\,
            I => \N__8090\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__8096\,
            I => \N__8087\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__8095\,
            I => \N__8084\
        );

    \I__1122\ : InMux
    port map (
            O => \N__8094\,
            I => \N__8077\
        );

    \I__1121\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8077\
        );

    \I__1120\ : Span4Mux_v
    port map (
            O => \N__8090\,
            I => \N__8074\
        );

    \I__1119\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8065\
        );

    \I__1118\ : InMux
    port map (
            O => \N__8084\,
            I => \N__8065\
        );

    \I__1117\ : InMux
    port map (
            O => \N__8083\,
            I => \N__8065\
        );

    \I__1116\ : InMux
    port map (
            O => \N__8082\,
            I => \N__8065\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__8077\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1114\ : Odrv4
    port map (
            O => \N__8074\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__8065\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__8058\,
            I => \N__8055\
        );

    \I__1111\ : InMux
    port map (
            O => \N__8055\,
            I => \N__8052\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__8052\,
            I => \N__8049\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__8049\,
            I => \uu2.mem0.w_addr_0\
        );

    \I__1108\ : InMux
    port map (
            O => \N__8046\,
            I => \N__8043\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__8043\,
            I => \N__8040\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__8040\,
            I => \uu2.r_data_wire_1\
        );

    \I__1105\ : InMux
    port map (
            O => \N__8037\,
            I => \N__8034\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__8034\,
            I => \N__8031\
        );

    \I__1103\ : Odrv4
    port map (
            O => \N__8031\,
            I => \uu2.r_data_wire_2\
        );

    \I__1102\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8025\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__8025\,
            I => \N__8022\
        );

    \I__1100\ : Span4Mux_v
    port map (
            O => \N__8022\,
            I => \N__8019\
        );

    \I__1099\ : Odrv4
    port map (
            O => \N__8019\,
            I => \uu2.r_data_wire_0\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__8016\,
            I => \uu2.mem0.N_7_0_cascade_\
        );

    \I__1097\ : InMux
    port map (
            O => \N__8013\,
            I => \N__8010\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__8010\,
            I => \uu2.mem0.w_data_1\
        );

    \I__1095\ : InMux
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__8004\,
            I => \N__8001\
        );

    \I__1093\ : Odrv4
    port map (
            O => \N__8001\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_22\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__7998\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_\
        );

    \I__1091\ : InMux
    port map (
            O => \N__7995\,
            I => \N__7992\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__7992\,
            I => \uu2.mem0.w_data_4\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1088\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7983\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__7983\,
            I => \uu2.mem0.G_14_0_a6_0_0_1\
        );

    \I__1086\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__7977\,
            I => \uu2.mem0.w_data_3\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__7974\,
            I => \uu2.N_326_0_cascade_\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__7971\,
            I => \uu2.vbuf_raddr.un469_ci_0_cascade_\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__7968\,
            I => \N__7965\
        );

    \I__1081\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7962\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__7962\,
            I => \N__7958\
        );

    \I__1079\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7955\
        );

    \I__1078\ : Odrv4
    port map (
            O => \N__7958\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__7955\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1075\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__7944\,
            I => \N__7941\
        );

    \I__1073\ : Span4Mux_h
    port map (
            O => \N__7941\,
            I => \N__7935\
        );

    \I__1072\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7932\
        );

    \I__1071\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7927\
        );

    \I__1070\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7927\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__7935\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__7932\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__7927\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__7920\,
            I => \N__7915\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__7919\,
            I => \N__7911\
        );

    \I__1064\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7908\
        );

    \I__1063\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7905\
        );

    \I__1062\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7899\
        );

    \I__1061\ : InMux
    port map (
            O => \N__7911\,
            I => \N__7899\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__7908\,
            I => \N__7894\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__7905\,
            I => \N__7894\
        );

    \I__1058\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7891\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__7899\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1056\ : Odrv4
    port map (
            O => \N__7894\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__7891\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1054\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7881\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__7881\,
            I => \uu2.vbuf_raddr.un447_ci_3\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__7878\,
            I => \N__7875\
        );

    \I__1051\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7872\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__7872\,
            I => \N__7866\
        );

    \I__1049\ : InMux
    port map (
            O => \N__7871\,
            I => \N__7863\
        );

    \I__1048\ : InMux
    port map (
            O => \N__7870\,
            I => \N__7858\
        );

    \I__1047\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7858\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__7866\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__7863\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__7858\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__7851\,
            I => \uu2.vbuf_raddr.un447_ci_3_cascade_\
        );

    \I__1042\ : InMux
    port map (
            O => \N__7848\,
            I => \N__7840\
        );

    \I__1041\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7840\
        );

    \I__1040\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7835\
        );

    \I__1039\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7835\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__7840\,
            I => \uu2.un425_ci_0\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__7835\,
            I => \uu2.un425_ci_0\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__7830\,
            I => \N__7827\
        );

    \I__1035\ : InMux
    port map (
            O => \N__7827\,
            I => \N__7824\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__7824\,
            I => \N__7819\
        );

    \I__1033\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7816\
        );

    \I__1032\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7813\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__7819\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__7816\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__7813\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__7806\,
            I => \N__7803\
        );

    \I__1027\ : InMux
    port map (
            O => \N__7803\,
            I => \N__7798\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__7802\,
            I => \N__7795\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__7801\,
            I => \N__7792\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__7798\,
            I => \N__7789\
        );

    \I__1023\ : InMux
    port map (
            O => \N__7795\,
            I => \N__7784\
        );

    \I__1022\ : InMux
    port map (
            O => \N__7792\,
            I => \N__7784\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__7789\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__7784\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1019\ : InMux
    port map (
            O => \N__7779\,
            I => \N__7776\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__7776\,
            I => \N__7773\
        );

    \I__1017\ : Odrv4
    port map (
            O => \N__7773\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_21\
        );

    \I__1016\ : InMux
    port map (
            O => \N__7770\,
            I => \N__7767\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__7767\,
            I => \uu2.mem0.w_data_0\
        );

    \I__1014\ : InMux
    port map (
            O => \N__7764\,
            I => \N__7761\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__7761\,
            I => \N__7758\
        );

    \I__1012\ : Span4Mux_v
    port map (
            O => \N__7758\,
            I => \N__7755\
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__7755\,
            I => \uu2.mem0.w_data_ns_1_5\
        );

    \I__1010\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7749\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__7749\,
            I => \uu2.mem0.w_data_5\
        );

    \I__1008\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7743\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__7743\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_17\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__7740\,
            I => \uu2.mem0.G_14_0_a6_0_cascade_\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__7737\,
            I => \N__7734\
        );

    \I__1004\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7730\
        );

    \I__1003\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7727\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__7730\,
            I => \N__7721\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__7727\,
            I => \N__7721\
        );

    \I__1000\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7717\
        );

    \I__999\ : Span4Mux_v
    port map (
            O => \N__7721\,
            I => \N__7714\
        );

    \I__998\ : InMux
    port map (
            O => \N__7720\,
            I => \N__7711\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__7717\,
            I => \Lab_UT.secuu0.un197_ci_9\
        );

    \I__996\ : Odrv4
    port map (
            O => \N__7714\,
            I => \Lab_UT.secuu0.un197_ci_9\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__7711\,
            I => \Lab_UT.secuu0.un197_ci_9\
        );

    \I__994\ : InMux
    port map (
            O => \N__7704\,
            I => \N__7699\
        );

    \I__993\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7696\
        );

    \I__992\ : InMux
    port map (
            O => \N__7702\,
            I => \N__7693\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__7699\,
            I => \N__7690\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__7696\,
            I => \Lab_UT.secuu0.l_countZ0Z_12\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__7693\,
            I => \Lab_UT.secuu0.l_countZ0Z_12\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__7690\,
            I => \Lab_UT.secuu0.l_countZ0Z_12\
        );

    \I__987\ : InMux
    port map (
            O => \N__7683\,
            I => \N__7677\
        );

    \I__986\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7677\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__7677\,
            I => \N__7667\
        );

    \I__984\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7662\
        );

    \I__983\ : InMux
    port map (
            O => \N__7675\,
            I => \N__7662\
        );

    \I__982\ : InMux
    port map (
            O => \N__7674\,
            I => \N__7659\
        );

    \I__981\ : InMux
    port map (
            O => \N__7673\,
            I => \N__7654\
        );

    \I__980\ : InMux
    port map (
            O => \N__7672\,
            I => \N__7654\
        );

    \I__979\ : InMux
    port map (
            O => \N__7671\,
            I => \N__7650\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__7670\,
            I => \N__7647\
        );

    \I__977\ : Span4Mux_v
    port map (
            O => \N__7667\,
            I => \N__7637\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__7662\,
            I => \N__7637\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__7659\,
            I => \N__7637\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__7654\,
            I => \N__7637\
        );

    \I__973\ : InMux
    port map (
            O => \N__7653\,
            I => \N__7634\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__7650\,
            I => \N__7631\
        );

    \I__971\ : InMux
    port map (
            O => \N__7647\,
            I => \N__7626\
        );

    \I__970\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7626\
        );

    \I__969\ : Span4Mux_h
    port map (
            O => \N__7637\,
            I => \N__7623\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__7634\,
            I => \N__7620\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__7631\,
            I => \Lab_UT.secuu0.un153_ci\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__7626\,
            I => \Lab_UT.secuu0.un153_ci\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__7623\,
            I => \Lab_UT.secuu0.un153_ci\
        );

    \I__964\ : Odrv12
    port map (
            O => \N__7620\,
            I => \Lab_UT.secuu0.un153_ci\
        );

    \I__963\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7608\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__7608\,
            I => \Lab_UT.secuu0.un208_ci_0\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__7605\,
            I => \N__7601\
        );

    \I__960\ : InMux
    port map (
            O => \N__7604\,
            I => \N__7598\
        );

    \I__959\ : InMux
    port map (
            O => \N__7601\,
            I => \N__7595\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__7598\,
            I => \N__7592\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__7595\,
            I => \Lab_UT.secuu0.l_countZ0Z_13\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__7592\,
            I => \Lab_UT.secuu0.l_countZ0Z_13\
        );

    \I__955\ : CEMux
    port map (
            O => \N__7587\,
            I => \N__7566\
        );

    \I__954\ : CEMux
    port map (
            O => \N__7586\,
            I => \N__7566\
        );

    \I__953\ : CEMux
    port map (
            O => \N__7585\,
            I => \N__7566\
        );

    \I__952\ : CEMux
    port map (
            O => \N__7584\,
            I => \N__7566\
        );

    \I__951\ : CEMux
    port map (
            O => \N__7583\,
            I => \N__7566\
        );

    \I__950\ : CEMux
    port map (
            O => \N__7582\,
            I => \N__7566\
        );

    \I__949\ : CEMux
    port map (
            O => \N__7581\,
            I => \N__7566\
        );

    \I__948\ : GlobalMux
    port map (
            O => \N__7566\,
            I => \N__7563\
        );

    \I__947\ : gio2CtrlBuf
    port map (
            O => \N__7563\,
            I => \Lab_UT.secuu0.un11_l_count_i_g\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__945\ : InMux
    port map (
            O => \N__7557\,
            I => \N__7546\
        );

    \I__944\ : InMux
    port map (
            O => \N__7556\,
            I => \N__7546\
        );

    \I__943\ : InMux
    port map (
            O => \N__7555\,
            I => \N__7546\
        );

    \I__942\ : InMux
    port map (
            O => \N__7554\,
            I => \N__7541\
        );

    \I__941\ : InMux
    port map (
            O => \N__7553\,
            I => \N__7541\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__7546\,
            I => \N__7535\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__7541\,
            I => \N__7535\
        );

    \I__938\ : InMux
    port map (
            O => \N__7540\,
            I => \N__7532\
        );

    \I__937\ : Span4Mux_h
    port map (
            O => \N__7535\,
            I => \N__7529\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__7532\,
            I => \Lab_UT.secuu0.l_precountZ0Z_0\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__7529\,
            I => \Lab_UT.secuu0.l_precountZ0Z_0\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__7524\,
            I => \uu2.un425_ci_0_cascade_\
        );

    \I__933\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7518\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__7518\,
            I => \N__7512\
        );

    \I__931\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7507\
        );

    \I__930\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7507\
        );

    \I__929\ : InMux
    port map (
            O => \N__7515\,
            I => \N__7504\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__7512\,
            I => \Lab_UT.secuu0.l_countZ0Z_10\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__7507\,
            I => \Lab_UT.secuu0.l_countZ0Z_10\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__7504\,
            I => \Lab_UT.secuu0.l_countZ0Z_10\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__7497\,
            I => \Lab_UT.secuu0.un186_ci_0_cascade_\
        );

    \I__924\ : InMux
    port map (
            O => \N__7494\,
            I => \N__7490\
        );

    \I__923\ : InMux
    port map (
            O => \N__7493\,
            I => \N__7485\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__7490\,
            I => \N__7480\
        );

    \I__921\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7477\
        );

    \I__920\ : InMux
    port map (
            O => \N__7488\,
            I => \N__7474\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__7485\,
            I => \N__7471\
        );

    \I__918\ : InMux
    port map (
            O => \N__7484\,
            I => \N__7466\
        );

    \I__917\ : InMux
    port map (
            O => \N__7483\,
            I => \N__7466\
        );

    \I__916\ : Span4Mux_s3_v
    port map (
            O => \N__7480\,
            I => \N__7457\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__7477\,
            I => \N__7457\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__7474\,
            I => \N__7457\
        );

    \I__913\ : Span4Mux_v
    port map (
            O => \N__7471\,
            I => \N__7457\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__7466\,
            I => \Lab_UT.secuu0.l_countZ0Z_8\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__7457\,
            I => \Lab_UT.secuu0.l_countZ0Z_8\
        );

    \I__910\ : InMux
    port map (
            O => \N__7452\,
            I => \N__7448\
        );

    \I__909\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7445\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__7448\,
            I => \N__7441\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__7445\,
            I => \N__7436\
        );

    \I__906\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7433\
        );

    \I__905\ : Span4Mux_h
    port map (
            O => \N__7441\,
            I => \N__7430\
        );

    \I__904\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7425\
        );

    \I__903\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7425\
        );

    \I__902\ : Span4Mux_h
    port map (
            O => \N__7436\,
            I => \N__7422\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__7433\,
            I => \Lab_UT.secuu0.l_countZ0Z_9\
        );

    \I__900\ : Odrv4
    port map (
            O => \N__7430\,
            I => \Lab_UT.secuu0.l_countZ0Z_9\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__7425\,
            I => \Lab_UT.secuu0.l_countZ0Z_9\
        );

    \I__898\ : Odrv4
    port map (
            O => \N__7422\,
            I => \Lab_UT.secuu0.l_countZ0Z_9\
        );

    \I__897\ : InMux
    port map (
            O => \N__7413\,
            I => \N__7408\
        );

    \I__896\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7403\
        );

    \I__895\ : InMux
    port map (
            O => \N__7411\,
            I => \N__7403\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__7408\,
            I => \N__7400\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__7403\,
            I => \Lab_UT.secuu0.l_countZ0Z_7\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__7400\,
            I => \Lab_UT.secuu0.l_countZ0Z_7\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__7395\,
            I => \N__7391\
        );

    \I__890\ : InMux
    port map (
            O => \N__7394\,
            I => \N__7387\
        );

    \I__889\ : InMux
    port map (
            O => \N__7391\,
            I => \N__7384\
        );

    \I__888\ : InMux
    port map (
            O => \N__7390\,
            I => \N__7381\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__7387\,
            I => \N__7378\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__7384\,
            I => \Lab_UT.secuu0.l_countZ0Z_3\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__7381\,
            I => \Lab_UT.secuu0.l_countZ0Z_3\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__7378\,
            I => \Lab_UT.secuu0.l_countZ0Z_3\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__7371\,
            I => \N__7368\
        );

    \I__882\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7364\
        );

    \I__881\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7360\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__7364\,
            I => \N__7357\
        );

    \I__879\ : InMux
    port map (
            O => \N__7363\,
            I => \N__7354\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__7360\,
            I => \Lab_UT.secuu0.l_countZ0Z_11\
        );

    \I__877\ : Odrv4
    port map (
            O => \N__7357\,
            I => \Lab_UT.secuu0.l_countZ0Z_11\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__7354\,
            I => \Lab_UT.secuu0.l_countZ0Z_11\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__7347\,
            I => \Lab_UT.secuu0.un4_l_count_11_cascade_\
        );

    \I__874\ : InMux
    port map (
            O => \N__7344\,
            I => \N__7338\
        );

    \I__873\ : InMux
    port map (
            O => \N__7343\,
            I => \N__7335\
        );

    \I__872\ : InMux
    port map (
            O => \N__7342\,
            I => \N__7330\
        );

    \I__871\ : InMux
    port map (
            O => \N__7341\,
            I => \N__7330\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__7338\,
            I => \N__7327\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__7335\,
            I => \Lab_UT.secuu0.l_countZ0Z_6\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__7330\,
            I => \Lab_UT.secuu0.l_countZ0Z_6\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__7327\,
            I => \Lab_UT.secuu0.l_countZ0Z_6\
        );

    \I__866\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7317\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__7317\,
            I => \N__7314\
        );

    \I__864\ : Odrv4
    port map (
            O => \N__7314\,
            I => \Lab_UT.secuu0.un4_l_count_16\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__7311\,
            I => \N__7307\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__7310\,
            I => \N__7303\
        );

    \I__861\ : InMux
    port map (
            O => \N__7307\,
            I => \N__7300\
        );

    \I__860\ : InMux
    port map (
            O => \N__7306\,
            I => \N__7295\
        );

    \I__859\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7295\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__7300\,
            I => \Lab_UT.secuu0.l_countZ0Z_17\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__7295\,
            I => \Lab_UT.secuu0.l_countZ0Z_17\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__7290\,
            I => \N__7285\
        );

    \I__855\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7282\
        );

    \I__854\ : InMux
    port map (
            O => \N__7288\,
            I => \N__7277\
        );

    \I__853\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7277\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__7282\,
            I => \N__7274\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__7277\,
            I => \N__7271\
        );

    \I__850\ : Span4Mux_h
    port map (
            O => \N__7274\,
            I => \N__7268\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__7271\,
            I => \Lab_UT.secuu0.un241_ci_2\
        );

    \I__848\ : Odrv4
    port map (
            O => \N__7268\,
            I => \Lab_UT.secuu0.un241_ci_2\
        );

    \I__847\ : InMux
    port map (
            O => \N__7263\,
            I => \N__7259\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__7262\,
            I => \N__7254\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__7259\,
            I => \N__7251\
        );

    \I__844\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7246\
        );

    \I__843\ : InMux
    port map (
            O => \N__7257\,
            I => \N__7246\
        );

    \I__842\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7243\
        );

    \I__841\ : Span4Mux_v
    port map (
            O => \N__7251\,
            I => \N__7240\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__7246\,
            I => \Lab_UT.secuu0.l_countZ0Z_16\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__7243\,
            I => \Lab_UT.secuu0.l_countZ0Z_16\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__7240\,
            I => \Lab_UT.secuu0.l_countZ0Z_16\
        );

    \I__837\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7230\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__7230\,
            I => \Lab_UT.secuu0.un263_ci\
        );

    \I__835\ : InMux
    port map (
            O => \N__7227\,
            I => \N__7223\
        );

    \I__834\ : InMux
    port map (
            O => \N__7226\,
            I => \N__7220\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__7223\,
            I => \Lab_UT.secuu0.l_countZ0Z_18\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__7220\,
            I => \Lab_UT.secuu0.l_countZ0Z_18\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__7215\,
            I => \uu2.un2_w_addr_user_5_cascade_\
        );

    \I__830\ : InMux
    port map (
            O => \N__7212\,
            I => \N__7209\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__7209\,
            I => \uu2.un2_w_addr_user_4\
        );

    \I__828\ : InMux
    port map (
            O => \N__7206\,
            I => \N__7203\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__7203\,
            I => \N__7200\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__7200\,
            I => \uu2.un2_w_addr_user\
        );

    \I__825\ : InMux
    port map (
            O => \N__7197\,
            I => \N__7180\
        );

    \I__824\ : InMux
    port map (
            O => \N__7196\,
            I => \N__7180\
        );

    \I__823\ : InMux
    port map (
            O => \N__7195\,
            I => \N__7180\
        );

    \I__822\ : InMux
    port map (
            O => \N__7194\,
            I => \N__7180\
        );

    \I__821\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7169\
        );

    \I__820\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7169\
        );

    \I__819\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7169\
        );

    \I__818\ : InMux
    port map (
            O => \N__7190\,
            I => \N__7169\
        );

    \I__817\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7169\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__7180\,
            I => \uu2.un27_w_addr_user_i\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__7169\,
            I => \uu2.un27_w_addr_user_i\
        );

    \I__814\ : SRMux
    port map (
            O => \N__7164\,
            I => \N__7161\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__7161\,
            I => \N__7157\
        );

    \I__812\ : SRMux
    port map (
            O => \N__7160\,
            I => \N__7154\
        );

    \I__811\ : Span4Mux_v
    port map (
            O => \N__7157\,
            I => \N__7151\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__7154\,
            I => \N__7148\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__7151\,
            I => \uu2.w_addr_user_RNIKHHELZ0Z_2\
        );

    \I__808\ : Odrv4
    port map (
            O => \N__7148\,
            I => \uu2.w_addr_user_RNIKHHELZ0Z_2\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__7143\,
            I => \N__7140\
        );

    \I__806\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7137\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__7137\,
            I => \uu2.o_adder_vbuf_w_addr_user_3\
        );

    \I__804\ : InMux
    port map (
            O => \N__7134\,
            I => \N__7124\
        );

    \I__803\ : InMux
    port map (
            O => \N__7133\,
            I => \N__7124\
        );

    \I__802\ : InMux
    port map (
            O => \N__7132\,
            I => \N__7121\
        );

    \I__801\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7118\
        );

    \I__800\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7115\
        );

    \I__799\ : InMux
    port map (
            O => \N__7129\,
            I => \N__7112\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__7124\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__7121\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__7118\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__7115\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__7112\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__7101\,
            I => \N__7096\
        );

    \I__792\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7089\
        );

    \I__791\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7089\
        );

    \I__790\ : InMux
    port map (
            O => \N__7096\,
            I => \N__7086\
        );

    \I__789\ : InMux
    port map (
            O => \N__7095\,
            I => \N__7083\
        );

    \I__788\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7080\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__7089\,
            I => \uu2.un425_ci\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__7086\,
            I => \uu2.un425_ci\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__7083\,
            I => \uu2.un425_ci\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__7080\,
            I => \uu2.un425_ci\
        );

    \I__783\ : InMux
    port map (
            O => \N__7071\,
            I => \N__7068\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__7068\,
            I => \N__7065\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__7065\,
            I => \uu2.r_data_wire_3\
        );

    \I__780\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7059\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__7059\,
            I => \uu2.un1_w_user_cr_5Z0Z_1\
        );

    \I__778\ : CascadeMux
    port map (
            O => \N__7056\,
            I => \Lab_UT_L3_tx_data_2_0_cascade_\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__7053\,
            I => \N__7049\
        );

    \I__776\ : InMux
    port map (
            O => \N__7052\,
            I => \N__7044\
        );

    \I__775\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7044\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__7044\,
            I => \uu2.un1_w_user_crZ0Z_5\
        );

    \I__773\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7038\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__7038\,
            I => \N__7034\
        );

    \I__771\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7031\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__7034\,
            I => \Lab_UT_L3_tx_data_0_6\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__7031\,
            I => \Lab_UT_L3_tx_data_0_6\
        );

    \I__768\ : InMux
    port map (
            O => \N__7026\,
            I => \N__7023\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__7023\,
            I => \uu2.mem0.w_data_6\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__7020\,
            I => \N__7016\
        );

    \I__765\ : InMux
    port map (
            O => \N__7019\,
            I => \N__7011\
        );

    \I__764\ : InMux
    port map (
            O => \N__7016\,
            I => \N__7008\
        );

    \I__763\ : InMux
    port map (
            O => \N__7015\,
            I => \N__7003\
        );

    \I__762\ : InMux
    port map (
            O => \N__7014\,
            I => \N__7003\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__7011\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__7008\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__7003\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__6996\,
            I => \N__6993\
        );

    \I__757\ : InMux
    port map (
            O => \N__6993\,
            I => \N__6990\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__6990\,
            I => \uu2.mem0.w_addr_8\
        );

    \I__755\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6984\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__6984\,
            I => \Lab_UT_L3_tx_data_2_0\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__6981\,
            I => \N__6978\
        );

    \I__752\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6975\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__6975\,
            I => \uu2.mem0.w_addr_1\
        );

    \I__750\ : InMux
    port map (
            O => \N__6972\,
            I => \N__6969\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__6969\,
            I => \N__6963\
        );

    \I__748\ : InMux
    port map (
            O => \N__6968\,
            I => \N__6958\
        );

    \I__747\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6958\
        );

    \I__746\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6955\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__6963\,
            I => \L3_tx_data_2\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__6958\,
            I => \L3_tx_data_2\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__6955\,
            I => \L3_tx_data_2\
        );

    \I__742\ : InMux
    port map (
            O => \N__6948\,
            I => \N__6945\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__6945\,
            I => \uu2.mem0.w_data_2\
        );

    \I__740\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6936\
        );

    \I__739\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6936\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__6936\,
            I => \uu2.un27_w_addr_user_0\
        );

    \I__737\ : InMux
    port map (
            O => \N__6933\,
            I => \N__6928\
        );

    \I__736\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6925\
        );

    \I__735\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6922\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__6928\,
            I => \Lab_UT.dspStr.cntZ0Z_0\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__6925\,
            I => \Lab_UT.dspStr.cntZ0Z_0\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__6922\,
            I => \Lab_UT.dspStr.cntZ0Z_0\
        );

    \I__731\ : InMux
    port map (
            O => \N__6915\,
            I => \N__6912\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__6912\,
            I => \uu2.un1_w_user_lfZ0Z_1\
        );

    \I__729\ : InMux
    port map (
            O => \N__6909\,
            I => \N__6906\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__6906\,
            I => \uu2.un1_w_user_lfZ0Z_3\
        );

    \I__727\ : InMux
    port map (
            O => \N__6903\,
            I => \N__6900\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__6900\,
            I => \uu2.un1_w_user_cr_0_0\
        );

    \I__725\ : InMux
    port map (
            O => \N__6897\,
            I => \N__6894\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__6894\,
            I => \uu2.un1_w_user_crZ0Z_2\
        );

    \I__723\ : InMux
    port map (
            O => \N__6891\,
            I => \N__6888\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__6888\,
            I => \L3_tx_data_rdy\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__6885\,
            I => \uu2.un1_w_user_crZ0Z_2_cascade_\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__6882\,
            I => \uu2.un19_w_addr_userZ0Z_0_cascade_\
        );

    \I__719\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6873\
        );

    \I__718\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6873\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__6873\,
            I => \L3_tx_data_7\
        );

    \I__716\ : InMux
    port map (
            O => \N__6870\,
            I => \N__6867\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__6867\,
            I => \N__6864\
        );

    \I__714\ : Span4Mux_h
    port map (
            O => \N__6864\,
            I => \N__6861\
        );

    \I__713\ : Odrv4
    port map (
            O => \N__6861\,
            I => \uu2.mem0.w_data_7\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__6858\,
            I => \Lab_UT.dspStr.cnt11_1_cascade_\
        );

    \I__711\ : InMux
    port map (
            O => \N__6855\,
            I => \N__6851\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__6854\,
            I => \N__6848\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__6851\,
            I => \N__6845\
        );

    \I__708\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6842\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__6845\,
            I => \Lab_UT.dspStr.cnt11_0_i\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__6842\,
            I => \Lab_UT.dspStr.cnt11_0_i\
        );

    \I__705\ : IoInMux
    port map (
            O => \N__6837\,
            I => \N__6834\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__6834\,
            I => \N__6831\
        );

    \I__703\ : IoSpan4Mux
    port map (
            O => \N__6831\,
            I => \N__6828\
        );

    \I__702\ : Span4Mux_s2_h
    port map (
            O => \N__6828\,
            I => \N__6825\
        );

    \I__701\ : Odrv4
    port map (
            O => \N__6825\,
            I => \Lab_UT.secuu0.un11_l_count_i\
        );

    \I__700\ : InMux
    port map (
            O => \N__6822\,
            I => \N__6819\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__6819\,
            I => \Lab_UT_dspStr_un29_dOut_0\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__6816\,
            I => \N__6811\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__6815\,
            I => \N__6808\
        );

    \I__696\ : InMux
    port map (
            O => \N__6814\,
            I => \N__6801\
        );

    \I__695\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6801\
        );

    \I__694\ : InMux
    port map (
            O => \N__6808\,
            I => \N__6801\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__6801\,
            I => \Lab_UT.secuu0.l_precountZ0Z_3\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__6798\,
            I => \N__6793\
        );

    \I__691\ : InMux
    port map (
            O => \N__6797\,
            I => \N__6785\
        );

    \I__690\ : InMux
    port map (
            O => \N__6796\,
            I => \N__6785\
        );

    \I__689\ : InMux
    port map (
            O => \N__6793\,
            I => \N__6785\
        );

    \I__688\ : InMux
    port map (
            O => \N__6792\,
            I => \N__6782\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__6785\,
            I => \Lab_UT.secuu0.l_countZ0Z_1\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__6782\,
            I => \Lab_UT.secuu0.l_countZ0Z_1\
        );

    \I__685\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6762\
        );

    \I__684\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6762\
        );

    \I__683\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6762\
        );

    \I__682\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6762\
        );

    \I__681\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6762\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__6762\,
            I => \Lab_UT.secuu0.l_precountZ0Z_1\
        );

    \I__679\ : InMux
    port map (
            O => \N__6759\,
            I => \N__6753\
        );

    \I__678\ : InMux
    port map (
            O => \N__6758\,
            I => \N__6748\
        );

    \I__677\ : InMux
    port map (
            O => \N__6757\,
            I => \N__6748\
        );

    \I__676\ : InMux
    port map (
            O => \N__6756\,
            I => \N__6745\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__6753\,
            I => \Lab_UT.secuu0.l_countZ0Z_2\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__6748\,
            I => \Lab_UT.secuu0.l_countZ0Z_2\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__6745\,
            I => \Lab_UT.secuu0.l_countZ0Z_2\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__6738\,
            I => \N__6732\
        );

    \I__671\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6723\
        );

    \I__670\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6723\
        );

    \I__669\ : InMux
    port map (
            O => \N__6735\,
            I => \N__6723\
        );

    \I__668\ : InMux
    port map (
            O => \N__6732\,
            I => \N__6723\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__6723\,
            I => \Lab_UT.secuu0.l_precountZ0Z_2\
        );

    \I__666\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6707\
        );

    \I__665\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6707\
        );

    \I__664\ : InMux
    port map (
            O => \N__6718\,
            I => \N__6707\
        );

    \I__663\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6707\
        );

    \I__662\ : InMux
    port map (
            O => \N__6716\,
            I => \N__6704\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__6707\,
            I => \Lab_UT.secuu0.l_countZ0Z_0\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__6704\,
            I => \Lab_UT.secuu0.l_countZ0Z_0\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__6699\,
            I => \Lab_UT.secuu0.un4_l_count_14_cascade_\
        );

    \I__658\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6691\
        );

    \I__657\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6686\
        );

    \I__656\ : InMux
    port map (
            O => \N__6694\,
            I => \N__6686\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__6691\,
            I => \N__6680\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__6686\,
            I => \N__6680\
        );

    \I__653\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6677\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__6680\,
            I => \Lab_UT.secuu0.un4_l_count_0_8\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__6677\,
            I => \Lab_UT.secuu0.un4_l_count_0_8\
        );

    \I__650\ : InMux
    port map (
            O => \N__6672\,
            I => \N__6669\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__6669\,
            I => \Lab_UT.secuu0.un4_l_count_12\
        );

    \I__648\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6663\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__6663\,
            I => \Lab_UT.secuu0.un4_l_count_13\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__6660\,
            I => \Lab_UT.secuu0.un4_l_count_18_cascade_\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__6657\,
            I => \N__6654\
        );

    \I__644\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6651\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__6651\,
            I => \N__6648\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__6648\,
            I => \Lab_UT.secuu0.un230_ci_1\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__6645\,
            I => \N__6639\
        );

    \I__640\ : InMux
    port map (
            O => \N__6644\,
            I => \N__6636\
        );

    \I__639\ : InMux
    port map (
            O => \N__6643\,
            I => \N__6633\
        );

    \I__638\ : InMux
    port map (
            O => \N__6642\,
            I => \N__6627\
        );

    \I__637\ : InMux
    port map (
            O => \N__6639\,
            I => \N__6627\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__6636\,
            I => \N__6624\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__6633\,
            I => \N__6621\
        );

    \I__634\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6618\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__6627\,
            I => \Lab_UT.secuu0.un109_ci\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__6624\,
            I => \Lab_UT.secuu0.un109_ci\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__6621\,
            I => \Lab_UT.secuu0.un109_ci\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__6618\,
            I => \Lab_UT.secuu0.un109_ci\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__6609\,
            I => \Lab_UT.secuu0.un197_ci_9_cascade_\
        );

    \I__628\ : InMux
    port map (
            O => \N__6606\,
            I => \N__6600\
        );

    \I__627\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6593\
        );

    \I__626\ : InMux
    port map (
            O => \N__6604\,
            I => \N__6593\
        );

    \I__625\ : InMux
    port map (
            O => \N__6603\,
            I => \N__6593\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__6600\,
            I => \Lab_UT.secuu0.l_countZ0Z_14\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__6593\,
            I => \Lab_UT.secuu0.l_countZ0Z_14\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__6588\,
            I => \N__6583\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__6587\,
            I => \N__6580\
        );

    \I__620\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6573\
        );

    \I__619\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6573\
        );

    \I__618\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6573\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__6573\,
            I => \Lab_UT.secuu0.l_countZ0Z_15\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__6570\,
            I => \N__6565\
        );

    \I__615\ : InMux
    port map (
            O => \N__6569\,
            I => \N__6561\
        );

    \I__614\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6558\
        );

    \I__613\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6553\
        );

    \I__612\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6553\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__6561\,
            I => \Lab_UT.secuu0.l_countZ0Z_4\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__6558\,
            I => \Lab_UT.secuu0.l_countZ0Z_4\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__6553\,
            I => \Lab_UT.secuu0.l_countZ0Z_4\
        );

    \I__608\ : InMux
    port map (
            O => \N__6546\,
            I => \N__6541\
        );

    \I__607\ : InMux
    port map (
            O => \N__6545\,
            I => \N__6538\
        );

    \I__606\ : InMux
    port map (
            O => \N__6544\,
            I => \N__6535\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__6541\,
            I => \N__6532\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__6538\,
            I => \Lab_UT.secuu0.l_countZ0Z_5\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__6535\,
            I => \Lab_UT.secuu0.l_countZ0Z_5\
        );

    \I__602\ : Odrv4
    port map (
            O => \N__6532\,
            I => \Lab_UT.secuu0.l_countZ0Z_5\
        );

    \I__601\ : InMux
    port map (
            O => \N__6525\,
            I => \N__6522\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__6522\,
            I => \uart_RXD\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__6519\,
            I => \uu2.un447_ci_3_cascade_\
        );

    \I__598\ : InMux
    port map (
            O => \N__6516\,
            I => \N__6513\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__6513\,
            I => \uu2.o_adder_vbuf_w_addr_user_7\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__6510\,
            I => \N__6507\
        );

    \I__595\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6504\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__6504\,
            I => \N__6501\
        );

    \I__593\ : Span4Mux_v
    port map (
            O => \N__6501\,
            I => \N__6498\
        );

    \I__592\ : Odrv4
    port map (
            O => \N__6498\,
            I => \uu2.mem0.w_addr_6\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__6495\,
            I => \N__6492\
        );

    \I__590\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__6489\,
            I => \N__6486\
        );

    \I__588\ : Span4Mux_h
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__587\ : Odrv4
    port map (
            O => \N__6483\,
            I => \uu2.mem0.w_addr_7\
        );

    \I__586\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6473\
        );

    \I__585\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6464\
        );

    \I__584\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6464\
        );

    \I__583\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6464\
        );

    \I__582\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6464\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__6473\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__6464\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__579\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6452\
        );

    \I__578\ : InMux
    port map (
            O => \N__6458\,
            I => \N__6447\
        );

    \I__577\ : InMux
    port map (
            O => \N__6457\,
            I => \N__6447\
        );

    \I__576\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6442\
        );

    \I__575\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6442\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__6452\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__6447\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__6442\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__6435\,
            I => \N__6432\
        );

    \I__570\ : InMux
    port map (
            O => \N__6432\,
            I => \N__6428\
        );

    \I__569\ : InMux
    port map (
            O => \N__6431\,
            I => \N__6425\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__6428\,
            I => \uu2.un447_ci_3\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__6425\,
            I => \uu2.un447_ci_3\
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__6420\,
            I => \uu2.vbuf_w_addr_user.un469_ci_0_cascade_\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__6417\,
            I => \N__6414\
        );

    \I__564\ : InMux
    port map (
            O => \N__6414\,
            I => \N__6411\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__6411\,
            I => \uu2.o_adder_vbuf_w_addr_user_8\
        );

    \I__562\ : InMux
    port map (
            O => \N__6408\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_2\
        );

    \I__561\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__6402\,
            I => \N__6399\
        );

    \I__559\ : Odrv4
    port map (
            O => \N__6399\,
            I => \uu2.un1_w_user_lfZ0Z_4\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__6396\,
            I => \L3_tx_data_0_cascade_\
        );

    \I__557\ : InMux
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__6390\,
            I => \uu2.un1_w_user_lf_0\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__6387\,
            I => \uu2.un1_w_user_lf_0_cascade_\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__6384\,
            I => \Lab_UT_L3_tx_data_0_4_cascade_\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__6381\,
            I => \Lab_UT_dspStr_un29_dOut_0_cascade_\
        );

    \I__552\ : InMux
    port map (
            O => \N__6378\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_0\
        );

    \I__551\ : InMux
    port map (
            O => \N__6375\,
            I => \Lab_UT.dspStr.un1_cnt_3_cry_1\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__6372\,
            I => \N__6369\
        );

    \I__549\ : InMux
    port map (
            O => \N__6369\,
            I => \N__6366\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__6366\,
            I => \Lab_UT.secuu0.un142_ci_0\
        );

    \I__547\ : CascadeMux
    port map (
            O => \N__6363\,
            I => \N__6359\
        );

    \I__546\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6354\
        );

    \I__545\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6354\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__6354\,
            I => \Lab_UT.secuu0.un131_ci_3\
        );

    \I__543\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6348\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__6348\,
            I => \Lab_UT.secuu0.un87_ci\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__6345\,
            I => \Lab_UT.secuu0.un87_ci_cascade_\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__6342\,
            I => \Lab_UT.secuu0.un131_ci_3_cascade_\
        );

    \I__539\ : IoInMux
    port map (
            O => \N__6339\,
            I => \N__6336\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__6336\,
            I => \N__6333\
        );

    \I__537\ : IoSpan4Mux
    port map (
            O => \N__6333\,
            I => \N__6330\
        );

    \I__536\ : Odrv4
    port map (
            O => \N__6330\,
            I => clk_in_c
        );

    \INVuu2.w_addr_displaying_0C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_0C_net\,
            I => \N__13494\
        );

    \INVuu2.w_addr_displaying_2_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_2_rep1C_net\,
            I => \N__13499\
        );

    \INVuu2.w_addr_displaying_0_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_0_rep1C_net\,
            I => \N__13504\
        );

    \INVuu2.w_addr_displaying_4_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_4_rep1C_net\,
            I => \N__13520\
        );

    \INVuu2.w_addr_displaying_fast_3C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_3C_net\,
            I => \N__13498\
        );

    \INVuu2.w_addr_displaying_6_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_6_rep1C_net\,
            I => \N__13503\
        );

    \INVuu2.w_addr_displaying_6C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_6C_net\,
            I => \N__13512\
        );

    \INVuu2.w_addr_displaying_2C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_2C_net\,
            I => \N__13484\
        );

    \INVuu2.w_addr_displaying_4C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_4C_net\,
            I => \N__13492\
        );

    \INVuu2.w_addr_displaying_fast_4C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_4C_net\,
            I => \N__13497\
        );

    \INVuu2.w_addr_displaying_5C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_5C_net\,
            I => \N__13483\
        );

    \INVuu2.w_addr_displaying_1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_1C_net\,
            I => \N__13491\
        );

    \INVuu2.w_addr_user_3C\ : INV
    port map (
            O => \INVuu2.w_addr_user_3C_net\,
            I => \N__13507\
        );

    \INVuu2.w_addr_user_4C\ : INV
    port map (
            O => \INVuu2.w_addr_user_4C_net\,
            I => \N__13515\
        );

    \IN_MUX_bfv_7_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_2_0_\
        );

    \IN_MUX_bfv_6_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_1_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_8_0_\
        );

    \latticehx1k_pll_inst.PLLOUTCORE_derived_clock_RNIALC1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8142\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \Lab_UT.secuu0.delay_line_RNILBAI7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6837\,
            GLOBALBUFFEROUTPUT => \Lab_UT.secuu0.un11_l_count_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \resetGen.rst_RNI4PQ1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10931\,
            GLOBALBUFFEROUTPUT => rst_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_5_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__6643\,
            in1 => \N__6545\,
            in2 => \_gnd_net_\,
            in3 => \N__6569\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13548\,
            ce => \N__7583\,
            sr => \N__15898\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_3_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6544\,
            in2 => \_gnd_net_\,
            in3 => \N__6568\,
            lcout => \Lab_UT.secuu0.un131_ci_3\,
            ltout => \Lab_UT.secuu0.un131_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_7__un142_ci_0_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6342\,
            in3 => \N__7343\,
            lcout => \Lab_UT.secuu0.un142_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_15__un230_ci_1_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6696\,
            in1 => \N__7726\,
            in2 => \_gnd_net_\,
            in3 => \N__6606\,
            lcout => \Lab_UT.secuu0.un230_ci_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_3_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__6351\,
            in1 => \N__6759\,
            in2 => \N__7395\,
            in3 => \N__11044\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13545\,
            ce => \N__7582\,
            sr => \N__15896\
        );

    \Lab_UT.secuu0.l_count_7_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__11043\,
            in1 => \N__6642\,
            in2 => \N__6372\,
            in3 => \N__7412\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13545\,
            ce => \N__7582\,
            sr => \N__15896\
        );

    \Lab_UT.secuu0.l_count_6_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__7342\,
            in1 => \N__6362\,
            in2 => \N__6645\,
            in3 => \N__11042\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13545\,
            ce => \N__7582\,
            sr => \N__15896\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_8_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6632\,
            in1 => \N__7341\,
            in2 => \N__6363\,
            in3 => \N__7411\,
            lcout => \Lab_UT.secuu0.un153_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_6_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6757\,
            in1 => \N__6717\,
            in2 => \N__6798\,
            in3 => \N__7390\,
            lcout => \Lab_UT.secuu0.un109_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_1_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__6720\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6797\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13541\,
            ce => \N__7581\,
            sr => \N__15895\
        );

    \Lab_UT.secuu0.l_count_0_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6719\,
            in2 => \_gnd_net_\,
            in3 => \N__11045\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13541\,
            ce => \N__7581\,
            sr => \N__15895\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_1_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6718\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6796\,
            lcout => \Lab_UT.secuu0.un87_ci\,
            ltout => \Lab_UT.secuu0.un87_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_2_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__6758\,
            in1 => \_gnd_net_\,
            in2 => \N__6345\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13541\,
            ce => \N__7581\,
            sr => \N__15895\
        );

    \Lab_UT.secuu0.l_count_RNIFM2M_13_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7604\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7704\,
            lcout => \Lab_UT.secuu0.un4_l_count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNIMHJI1_2_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011111100111"
        )
    port map (
            in0 => \N__8562\,
            in1 => \N__8728\,
            in2 => \N__8666\,
            in3 => \N__8842\,
            lcout => OPEN,
            ltout => \Lab_UT_L3_tx_data_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_4_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6384\,
            in3 => \N__6966\,
            lcout => \uu2.un1_w_user_lfZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNIKFJI1_2_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110100001"
        )
    port map (
            in0 => \N__8561\,
            in1 => \N__8726\,
            in2 => \N__8665\,
            in3 => \N__10297\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.Lab3U00.q_esr_2_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9666\,
            lcout => \Lab_UT.rx_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13533\,
            ce => \N__9090\,
            sr => \N__15873\
        );

    \Lab_UT.dspStr.cnt_RNI57RQ_2_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8642\,
            in2 => \_gnd_net_\,
            in3 => \N__8560\,
            lcout => \Lab_UT_dspStr_un29_dOut_0\,
            ltout => \Lab_UT_dspStr_un29_dOut_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_0_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101111111"
        )
    port map (
            in0 => \N__8841\,
            in1 => \N__8727\,
            in2 => \N__6381\,
            in3 => \N__8774\,
            lcout => \uu2.un1_w_user_cr_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_0_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6932\,
            in2 => \N__6854\,
            in3 => \N__6855\,
            lcout => \Lab_UT.dspStr.cntZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => \Lab_UT.dspStr.un1_cnt_3_cry_0\,
            clk => \N__13528\,
            ce => 'H',
            sr => \N__15872\
        );

    \Lab_UT.dspStr.cnt_1_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8742\,
            in2 => \_gnd_net_\,
            in3 => \N__6378\,
            lcout => \Lab_UT_dspStr_cnt_1\,
            ltout => OPEN,
            carryin => \Lab_UT.dspStr.un1_cnt_3_cry_0\,
            carryout => \Lab_UT.dspStr.un1_cnt_3_cry_1\,
            clk => \N__13528\,
            ce => 'H',
            sr => \N__15872\
        );

    \Lab_UT.dspStr.cnt_2_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8574\,
            in2 => \_gnd_net_\,
            in3 => \N__6375\,
            lcout => \Lab_UT_dspStr_cnt_2\,
            ltout => OPEN,
            carryin => \Lab_UT.dspStr.un1_cnt_3_cry_1\,
            carryout => \Lab_UT.dspStr.un1_cnt_3_cry_2\,
            clk => \N__13528\,
            ce => 'H',
            sr => \N__15872\
        );

    \Lab_UT.dspStr.cnt_3_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8664\,
            in2 => \_gnd_net_\,
            in3 => \N__6408\,
            lcout => \Lab_UT_dspStr_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13528\,
            ce => 'H',
            sr => \N__15872\
        );

    \uu2.w_addr_user_RNIKHHEL_2_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__10938\,
            in1 => \N__6942\,
            in2 => \_gnd_net_\,
            in3 => \N__6393\,
            lcout => \uu2.w_addr_user_RNIKHHELZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNIIDJI1_0_2_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010100010"
        )
    port map (
            in0 => \N__8741\,
            in1 => \N__8660\,
            in2 => \N__10370\,
            in3 => \N__8570\,
            lcout => OPEN,
            ltout => \L3_tx_data_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8162\,
            in1 => \N__6405\,
            in2 => \N__6396\,
            in3 => \N__6909\,
            lcout => \uu2.un1_w_user_lf_0\,
            ltout => \uu2.un1_w_user_lf_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNILJEE01_2_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6941\,
            in2 => \N__6387\,
            in3 => \N__12399\,
            lcout => \uu2.un27_w_addr_user_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_4_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__7099\,
            in1 => \N__9371\,
            in2 => \_gnd_net_\,
            in3 => \N__7194\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_4C_net\,
            ce => 'H',
            sr => \N__7160\
        );

    \uu2.w_addr_user_8_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__7196\,
            in1 => \_gnd_net_\,
            in2 => \N__6417\,
            in3 => \N__7019\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_4C_net\,
            ce => 'H',
            sr => \N__7160\
        );

    \uu2.w_addr_user_7_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6516\,
            in1 => \N__6459\,
            in2 => \_gnd_net_\,
            in3 => \N__7195\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_4C_net\,
            ce => 'H',
            sr => \N__7160\
        );

    \uu2.w_addr_user_6_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__7197\,
            in1 => \N__7100\,
            in2 => \N__6435\,
            in3 => \N__6480\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_4C_net\,
            ce => 'H',
            sr => \N__7160\
        );

    \buart.Z_rx.hh_0_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6525\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_6__un447_ci_3_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__9322\,
            in1 => \N__9370\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.un447_ci_3\,
            ltout => \uu2.un447_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.result_1_7_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__6479\,
            in1 => \N__7094\,
            in2 => \N__6519\,
            in3 => \N__6458\,
            lcout => \uu2.o_adder_vbuf_w_addr_user_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12460\,
            in1 => \N__6477\,
            in2 => \_gnd_net_\,
            in3 => \N__12231\,
            lcout => \uu2.mem0.w_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6456\,
            in1 => \N__12461\,
            in2 => \_gnd_net_\,
            in3 => \N__16290\,
            lcout => \uu2.mem0.w_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIOGH7_8_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__7014\,
            in1 => \N__6455\,
            in2 => \_gnd_net_\,
            in3 => \N__6476\,
            lcout => \uu2.un2_w_addr_user_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_8__un469_ci_0_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6478\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6457\,
            lcout => OPEN,
            ltout => \uu2.vbuf_w_addr_user.un469_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.result_1_8_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__7015\,
            in1 => \N__6431\,
            in2 => \N__6420\,
            in3 => \N__7095\,
            lcout => \uu2.o_adder_vbuf_w_addr_user_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_9_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__7671\,
            in1 => \N__7494\,
            in2 => \_gnd_net_\,
            in3 => \N__7444\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13547\,
            ce => \N__7586\,
            sr => \N__15901\
        );

    \Lab_UT.secuu0.l_count_10_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__7440\,
            in1 => \N__7517\,
            in2 => \N__7670\,
            in3 => \N__7489\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13546\,
            ce => \N__7584\,
            sr => \N__15899\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_16__un241_ci_2_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6604\,
            in1 => \N__7720\,
            in2 => \N__6588\,
            in3 => \N__6694\,
            lcout => \Lab_UT.secuu0.un241_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_15_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__6586\,
            in1 => \N__7646\,
            in2 => \N__6657\,
            in3 => \N__11040\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13546\,
            ce => \N__7584\,
            sr => \N__15899\
        );

    \Lab_UT.secuu0.l_count_4_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__11041\,
            in1 => \_gnd_net_\,
            in2 => \N__6570\,
            in3 => \N__6644\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13546\,
            ce => \N__7584\,
            sr => \N__15899\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_12__un197_ci_9_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7516\,
            in1 => \N__7439\,
            in2 => \N__7371\,
            in3 => \N__7488\,
            lcout => \Lab_UT.secuu0.un197_ci_9\,
            ltout => \Lab_UT.secuu0.un197_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_14_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__6695\,
            in1 => \N__7674\,
            in2 => \N__6609\,
            in3 => \N__6605\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13546\,
            ce => \N__7584\,
            sr => \N__15899\
        );

    \Lab_UT.secuu0.l_count_RNIGLN81_15_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6603\,
            in1 => \N__7515\,
            in2 => \N__6587\,
            in3 => \N__6564\,
            lcout => \Lab_UT.secuu0.un4_l_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.delay_line_0_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6774\,
            in1 => \N__7555\,
            in2 => \N__6816\,
            in3 => \N__6735\,
            lcout => \Lab_UT.secuu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13542\,
            ce => 'H',
            sr => \N__15897\
        );

    \Lab_UT.secuu0.l_precount_3_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__6737\,
            in1 => \N__6814\,
            in2 => \N__7560\,
            in3 => \N__6777\,
            lcout => \Lab_UT.secuu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13542\,
            ce => 'H',
            sr => \N__15897\
        );

    \Lab_UT.secuu0.l_count_RNI8TM21_5_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6773\,
            in1 => \N__6546\,
            in2 => \N__6815\,
            in3 => \N__6792\,
            lcout => \Lab_UT.secuu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_precount_1_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7554\,
            in2 => \_gnd_net_\,
            in3 => \N__6775\,
            lcout => \Lab_UT.secuu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13542\,
            ce => 'H',
            sr => \N__15897\
        );

    \Lab_UT.secuu0.l_precount_2_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__6776\,
            in1 => \N__7556\,
            in2 => \_gnd_net_\,
            in3 => \N__6736\,
            lcout => \Lab_UT.secuu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13542\,
            ce => 'H',
            sr => \N__15897\
        );

    \Lab_UT.secuu0.l_count_RNI3II01_2_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7493\,
            in1 => \N__6756\,
            in2 => \N__6738\,
            in3 => \N__6716\,
            lcout => OPEN,
            ltout => \Lab_UT.secuu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_RNIOIEB2_16_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7553\,
            in1 => \N__7263\,
            in2 => \N__6699\,
            in3 => \N__6685\,
            lcout => OPEN,
            ltout => \Lab_UT.secuu0.un4_l_count_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_RNI82GM6_5_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6672\,
            in1 => \N__6666\,
            in2 => \N__6660\,
            in3 => \N__7320\,
            lcout => \Lab_UT.secuu0.un4_l_count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.Lab3U00.q_esr_0_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13599\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.rx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13534\,
            ce => \N__9083\,
            sr => \N__15875\
        );

    \Lab_UT.Lab3U00.q_esr_3_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9618\,
            lcout => \Lab_UT_rx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13534\,
            ce => \N__9083\,
            sr => \N__15875\
        );

    \Lab_UT.Lab3U00.q_esr_5_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8499\,
            lcout => \Lab_UT_rx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13534\,
            ce => \N__9083\,
            sr => \N__15875\
        );

    \Lab_UT.Lab3U00.q_esr_6_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9690\,
            lcout => \Lab_UT_rx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13534\,
            ce => \N__9083\,
            sr => \N__15875\
        );

    \Lab_UT.Lab3U00.q_esr_7_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9717\,
            lcout => \Lab_UT_rx_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13534\,
            ce => \N__9083\,
            sr => \N__15875\
        );

    \Lab_UT.Lab3U00.q_esr_4_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9642\,
            lcout => \Lab_UT_rx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13534\,
            ce => \N__9083\,
            sr => \N__15875\
        );

    \Lab_UT.dspStr.cnt_RNI11B71_2_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__16546\,
            in1 => \N__8654\,
            in2 => \N__13344\,
            in3 => \N__8565\,
            lcout => OPEN,
            ltout => \Lab_UT.dspStr.cnt11_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNI24622_0_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6931\,
            in2 => \N__6858\,
            in3 => \N__8724\,
            lcout => \Lab_UT.dspStr.cnt11_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.delay_line_RNILBAI7_1_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__10974\,
            in1 => \N__10988\,
            in2 => \_gnd_net_\,
            in3 => \N__11052\,
            lcout => \Lab_UT.secuu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_1_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__8772\,
            in1 => \N__8723\,
            in2 => \N__10225\,
            in3 => \N__6822\,
            lcout => \uu2.un1_w_user_lfZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_26_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110000100100"
        )
    port map (
            in0 => \N__8725\,
            in1 => \N__8653\,
            in2 => \N__8577\,
            in3 => \N__8773\,
            lcout => \uu2.mem0.w_data_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNIOJJI1_2_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110001000"
        )
    port map (
            in0 => \N__8563\,
            in1 => \N__8722\,
            in2 => \N__10155\,
            in3 => \N__8657\,
            lcout => \Lab_UT_L3_tx_data_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNIPKJI1_2_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8721\,
            in1 => \N__8652\,
            in2 => \N__10224\,
            in3 => \N__8564\,
            lcout => \L3_tx_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNILGJI1_2_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001111"
        )
    port map (
            in0 => \N__8650\,
            in1 => \N__8808\,
            in2 => \N__8745\,
            in3 => \N__8569\,
            lcout => \L3_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIG1C8B_2_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__6968\,
            in1 => \N__7206\,
            in2 => \N__7053\,
            in3 => \N__6897\,
            lcout => \uu2.un27_w_addr_user_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.rdy_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6933\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13522\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_5_1_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000110011"
        )
    port map (
            in0 => \N__10197\,
            in1 => \N__8737\,
            in2 => \N__8815\,
            in3 => \N__8649\,
            lcout => \uu2.un1_w_user_cr_5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_3_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8651\,
            in1 => \N__8754\,
            in2 => \N__10163\,
            in3 => \N__6915\,
            lcout => \uu2.un1_w_user_lfZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_2_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7037\,
            in1 => \N__6878\,
            in2 => \_gnd_net_\,
            in3 => \N__6903\,
            lcout => \uu2.un1_w_user_crZ0Z_2\,
            ltout => \uu2.un1_w_user_crZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un19_w_addr_user_0_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__6891\,
            in1 => \N__7052\,
            in2 => \N__6885\,
            in3 => \N__6967\,
            lcout => \uu2.un19_w_addr_userZ0Z_0\,
            ltout => \uu2.un19_w_addr_userZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_15_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6882\,
            in3 => \N__6879\,
            lcout => \uu2.mem0.w_data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dspStr.cnt_RNIIDJI1_2_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110011"
        )
    port map (
            in0 => \N__8729\,
            in1 => \N__8655\,
            in2 => \N__10369\,
            in3 => \N__8566\,
            lcout => \Lab_UT_L3_tx_data_2_0\,
            ltout => \Lab_UT_L3_tx_data_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_5_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__8567\,
            in1 => \N__7062\,
            in2 => \N__7056\,
            in3 => \N__8658\,
            lcout => \uu2.un1_w_user_crZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__7041\,
            in1 => \N__8927\,
            in2 => \_gnd_net_\,
            in3 => \N__12425\,
            lcout => \uu2.mem0.w_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12420\,
            in2 => \N__7020\,
            in3 => \N__12576\,
            lcout => \uu2.mem0.w_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_21_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8731\,
            in1 => \N__6987\,
            in2 => \_gnd_net_\,
            in3 => \N__8656\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_22_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000110001000"
        )
    port map (
            in0 => \N__8568\,
            in1 => \N__8730\,
            in2 => \N__8859\,
            in3 => \N__8659\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__7130\,
            in1 => \_gnd_net_\,
            in2 => \N__12462\,
            in3 => \N__14998\,
            lcout => \uu2.mem0.w_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12424\,
            in2 => \_gnd_net_\,
            in3 => \N__6972\,
            lcout => \uu2.mem0.w_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_3_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__8988\,
            in1 => \_gnd_net_\,
            in2 => \N__7143\,
            in3 => \N__7191\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_3C_net\,
            ce => 'H',
            sr => \N__7164\
        );

    \uu2.w_addr_user_1_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__7190\,
            in1 => \_gnd_net_\,
            in2 => \N__8095\,
            in3 => \N__7133\,
            lcout => \uu2.w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_3C_net\,
            ce => 'H',
            sr => \N__7164\
        );

    \uu2.w_addr_user_RNIDD1A_5_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8987\,
            in1 => \N__7129\,
            in2 => \N__9323\,
            in3 => \N__8082\,
            lcout => OPEN,
            ltout => \uu2.un2_w_addr_user_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIDMJM_2_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9365\,
            in1 => \N__9035\,
            in2 => \N__7215\,
            in3 => \N__7212\,
            lcout => \uu2.un2_w_addr_user\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_0_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8083\,
            in2 => \_gnd_net_\,
            in3 => \N__7189\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_3C_net\,
            ce => 'H',
            sr => \N__7164\
        );

    \uu2.w_addr_user_2_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__7192\,
            in1 => \N__9036\,
            in2 => \N__8096\,
            in3 => \N__7134\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_3C_net\,
            ce => 'H',
            sr => \N__7164\
        );

    \uu2.w_addr_user_5_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__9318\,
            in1 => \N__9366\,
            in2 => \N__7101\,
            in3 => \N__7193\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_3C_net\,
            ce => 'H',
            sr => \N__7164\
        );

    \uu2.vbuf_w_addr_user.result_1_3_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8094\,
            in1 => \N__8990\,
            in2 => \N__9047\,
            in3 => \N__7132\,
            lcout => \uu2.o_adder_vbuf_w_addr_user_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_4__un425_ci_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8989\,
            in1 => \N__7131\,
            in2 => \N__9046\,
            in3 => \N__8093\,
            lcout => \uu2.un425_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_esr_3_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7071\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13496\,
            ce => \N__11352\,
            sr => \N__15878\
        );

    \Lab_UT.secuu0.l_count_17_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__7258\,
            in1 => \N__7673\,
            in2 => \N__7311\,
            in3 => \N__7288\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13535\,
            ce => \N__7587\,
            sr => \N__15902\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_11__un186_ci_0_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7521\,
            in1 => \N__7483\,
            in2 => \_gnd_net_\,
            in3 => \N__7452\,
            lcout => OPEN,
            ltout => \Lab_UT.secuu0.un186_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_11_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__7675\,
            in1 => \N__7367\,
            in2 => \N__7497\,
            in3 => \N__11068\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13535\,
            ce => \N__7587\,
            sr => \N__15902\
        );

    \Lab_UT.secuu0.l_count_16_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__11069\,
            in1 => \N__7676\,
            in2 => \N__7290\,
            in3 => \N__7257\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13535\,
            ce => \N__7587\,
            sr => \N__15902\
        );

    \Lab_UT.secuu0.l_count_8_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7484\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7672\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13535\,
            ce => \N__7587\,
            sr => \N__15902\
        );

    \Lab_UT.secuu0.l_count_RNIRDS11_3_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__7451\,
            in1 => \N__7413\,
            in2 => \N__7310\,
            in3 => \N__7394\,
            lcout => OPEN,
            ltout => \Lab_UT.secuu0.un4_l_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_RNIOSIV1_18_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7226\,
            in1 => \N__7363\,
            in2 => \N__7347\,
            in3 => \N__7344\,
            lcout => \Lab_UT.secuu0.un4_l_count_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_13__un208_ci_0_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7733\,
            in2 => \_gnd_net_\,
            in3 => \N__7702\,
            lcout => \Lab_UT.secuu0.un208_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_18__un263_ci_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7306\,
            in1 => \N__7289\,
            in2 => \N__7262\,
            in3 => \N__7653\,
            lcout => \Lab_UT.secuu0.un263_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.l_count_18_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7233\,
            in1 => \N__7227\,
            in2 => \_gnd_net_\,
            in3 => \N__11072\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13523\,
            ce => \N__7585\,
            sr => \N__15900\
        );

    \Lab_UT.secuu0.l_count_12_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__7682\,
            in1 => \N__7703\,
            in2 => \N__7737\,
            in3 => \N__11070\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13523\,
            ce => \N__7585\,
            sr => \N__15900\
        );

    \Lab_UT.secuu0.l_count_13_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__11071\,
            in1 => \N__7683\,
            in2 => \N__7605\,
            in3 => \N__7611\,
            lcout => \Lab_UT.secuu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13523\,
            ce => \N__7585\,
            sr => \N__15900\
        );

    \Lab_UT.secuu0.l_precount_0_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7540\,
            lcout => \Lab_UT.secuu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13516\,
            ce => 'H',
            sr => \N__15877\
        );

    \uu2.r_addr_5_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__7848\,
            in1 => \N__7940\,
            in2 => \N__7919\,
            in3 => \N__11192\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13516\,
            ce => 'H',
            sr => \N__15877\
        );

    \uu2.r_addr_4_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__11191\,
            in1 => \N__7847\,
            in2 => \_gnd_net_\,
            in3 => \N__7914\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13516\,
            ce => 'H',
            sr => \N__15877\
        );

    \uu2.r_addr_0_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11255\,
            in2 => \_gnd_net_\,
            in3 => \N__11190\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13516\,
            ce => 'H',
            sr => \N__15877\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un425_ci_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11104\,
            in1 => \N__11314\,
            in2 => \N__7801\,
            in3 => \N__11253\,
            lcout => \uu2.un425_ci_0\,
            ltout => \uu2.un425_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_6_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__7939\,
            in1 => \N__7918\,
            in2 => \N__7524\,
            in3 => \N__7871\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13510\,
            ce => \N__11341\,
            sr => \N__15874\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un469_ci_0_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7822\,
            in2 => \_gnd_net_\,
            in3 => \N__7869\,
            lcout => OPEN,
            ltout => \uu2.vbuf_raddr.un469_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_8_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__7961\,
            in1 => \N__7884\,
            in2 => \N__7971\,
            in3 => \N__7845\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13510\,
            ce => \N__11341\,
            sr => \N__15874\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un447_ci_3_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7938\,
            in2 => \_gnd_net_\,
            in3 => \N__7904\,
            lcout => \uu2.vbuf_raddr.un447_ci_3\,
            ltout => \uu2.vbuf_raddr.un447_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_7_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__7870\,
            in1 => \N__7823\,
            in2 => \N__7851\,
            in3 => \N__7846\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13510\,
            ce => \N__11341\,
            sr => \N__15874\
        );

    \uu2.r_addr_esr_3_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11105\,
            in1 => \N__11315\,
            in2 => \N__7802\,
            in3 => \N__11254\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13510\,
            ce => \N__11341\,
            sr => \N__15874\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12476\,
            in1 => \N__7779\,
            in2 => \_gnd_net_\,
            in3 => \N__7746\,
            lcout => \uu2.mem0.w_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000011"
        )
    port map (
            in0 => \N__7764\,
            in1 => \N__9235\,
            in2 => \N__8931\,
            in3 => \N__12478\,
            lcout => \uu2.mem0.w_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_17_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__8918\,
            in1 => \_gnd_net_\,
            in2 => \N__9236\,
            in3 => \N__16202\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_37_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110011"
        )
    port map (
            in0 => \N__11439\,
            in1 => \N__12475\,
            in2 => \N__7989\,
            in3 => \N__8181\,
            lcout => OPEN,
            ltout => \uu2.mem0.G_14_0_a6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_24_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__10419\,
            in1 => \N__10560\,
            in2 => \N__7740\,
            in3 => \N__9096\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__11748\,
            in1 => \N__8940\,
            in2 => \N__8016\,
            in3 => \N__9249\,
            lcout => \uu2.mem0.w_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_18_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__8919\,
            in1 => \_gnd_net_\,
            in2 => \N__9237\,
            in3 => \N__16203\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8007\,
            in2 => \N__7998\,
            in3 => \N__12477\,
            lcout => \uu2.mem0.w_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNII1IB1_5_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000010000"
        )
    port map (
            in0 => \N__12229\,
            in1 => \N__12562\,
            in2 => \N__12322\,
            in3 => \N__16287\,
            lcout => \uu2.bitmap_pmux_1_1_a8_1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_49_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16288\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12563\,
            lcout => \uu2.mem0.G_14_0_a6_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101011111"
        )
    port map (
            in0 => \N__8151\,
            in1 => \N__9135\,
            in2 => \N__12482\,
            in3 => \N__9108\,
            lcout => \uu2.mem0.w_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI979P_3_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111011"
        )
    port map (
            in0 => \N__13083\,
            in1 => \N__14832\,
            in2 => \N__14987\,
            in3 => \N__14313\,
            lcout => \uu2.N_326_0\,
            ltout => \uu2.N_326_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0QUP1_6_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__12230\,
            in1 => \N__12561\,
            in2 => \N__7974\,
            in3 => \N__16286\,
            lcout => \uu2.bitmap_pmux_1_1_a8_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI28SI1_7_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__13856\,
            in1 => \N__14010\,
            in2 => \N__13035\,
            in3 => \N__14253\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_1_1_a8_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNITAMH5_7_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__8202\,
            in1 => \N__8196\,
            in2 => \N__8190\,
            in3 => \N__8187\,
            lcout => \uu2.bitmap_pmux_1_1_1_tz\,
            ltout => \uu2.bitmap_pmux_1_1_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_29_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010010000"
        )
    port map (
            in0 => \N__16289\,
            in1 => \N__12564\,
            in2 => \N__8175\,
            in3 => \N__11435\,
            lcout => \uu2.mem0.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_25_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100010001"
        )
    port map (
            in0 => \N__9217\,
            in1 => \N__8926\,
            in2 => \N__8172\,
            in3 => \N__12466\,
            lcout => \uu2.mem0.w_data_1_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_wr_en_0_i_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__8141\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12467\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12468\,
            in1 => \N__8100\,
            in2 => \_gnd_net_\,
            in3 => \N__16200\,
            lcout => \uu2.mem0.w_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__16098\,
            in1 => \N__16201\,
            in2 => \_gnd_net_\,
            in3 => \N__14961\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1C_net\,
            ce => 'H',
            sr => \N__15848\
        );

    \uu2.r_data_reg_esr_1_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8046\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13489\,
            ce => \N__11348\,
            sr => \N__15881\
        );

    \uu2.r_data_reg_esr_2_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8037\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13489\,
            ce => \N__11348\,
            sr => \N__15881\
        );

    \uu2.r_data_reg_esr_0_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8028\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13489\,
            ce => \N__11348\,
            sr => \N__15881\
        );

    \uu2.r_data_reg_esr_4_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8289\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13489\,
            ce => \N__11348\,
            sr => \N__15881\
        );

    \uu2.r_data_reg_esr_5_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8280\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13489\,
            ce => \N__11348\,
            sr => \N__15881\
        );

    \uu2.r_data_reg_esr_6_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13489\,
            ce => \N__11348\,
            sr => \N__15881\
        );

    \uu2.r_data_reg_esr_7_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8262\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13489\,
            ce => \N__11348\,
            sr => \N__15881\
        );

    \buart.Z_tx.shifter_1_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__11223\,
            in1 => \_gnd_net_\,
            in2 => \N__8253\,
            in3 => \N__8214\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13486\,
            ce => \N__9570\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_0_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8244\,
            in2 => \_gnd_net_\,
            in3 => \N__11221\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13486\,
            ce => \N__9570\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.uart_tx_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11222\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8238\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13486\,
            ce => \N__9570\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_2_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8220\,
            in1 => \N__8346\,
            in2 => \_gnd_net_\,
            in3 => \N__11224\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13486\,
            ce => \N__9570\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_3_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11225\,
            in1 => \N__8208\,
            in2 => \_gnd_net_\,
            in3 => \N__8328\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13486\,
            ce => \N__9570\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_4_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8340\,
            in1 => \N__8316\,
            in2 => \_gnd_net_\,
            in3 => \N__11226\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13486\,
            ce => \N__9570\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_5_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11227\,
            in1 => \N__8322\,
            in2 => \_gnd_net_\,
            in3 => \N__8304\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13486\,
            ce => \N__9570\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_6_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9159\,
            in1 => \N__8310\,
            in2 => \_gnd_net_\,
            in3 => \N__11228\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13486\,
            ce => \N__9570\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10105\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8405\,
            in2 => \_gnd_net_\,
            in3 => \N__8298\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10069\,
            in2 => \_gnd_net_\,
            in3 => \N__8295\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10013\,
            in2 => \_gnd_net_\,
            in3 => \N__8292\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_4_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101101001110"
        )
    port map (
            in0 => \N__8885\,
            in1 => \N__8427\,
            in2 => \N__9897\,
            in3 => \N__8433\,
            lcout => \buart__rx_bitcount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13536\,
            ce => \N__9825\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNI2B26_4_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8404\,
            in1 => \N__10070\,
            in2 => \N__10023\,
            in3 => \N__8426\,
            lcout => OPEN,
            ltout => \buart.Z_rx.N_144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNIBJOC_0_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9930\,
            in2 => \N__8430\,
            in3 => \N__10111\,
            lcout => \buart.Z_rx.N_41_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_i_0_o2_4_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__8425\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8403\,
            lcout => \N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_1_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101101001110"
        )
    port map (
            in0 => \N__8880\,
            in1 => \N__8412\,
            in2 => \N__9888\,
            in3 => \N__8406\,
            lcout => \buart__rx_bitcount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13529\,
            ce => \N__9824\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_2_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101011010"
        )
    port map (
            in0 => \N__10071\,
            in1 => \N__9875\,
            in2 => \N__8385\,
            in3 => \N__8881\,
            lcout => \buart__rx_bitcount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13529\,
            ce => \N__9824\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_3_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101011100"
        )
    port map (
            in0 => \N__9873\,
            in1 => \N__8376\,
            in2 => \N__8886\,
            in3 => \N__10014\,
            lcout => \buart__rx_bitcount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13529\,
            ce => \N__9824\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_0_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001101011010"
        )
    port map (
            in0 => \N__10112\,
            in1 => \N__9874\,
            in2 => \N__8369\,
            in3 => \N__8879\,
            lcout => \buart__rx_bitcount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13529\,
            ce => \N__9824\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_4_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8492\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13524\,
            ce => \N__13570\,
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_i_0_a3_5_4_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8491\,
            in1 => \N__9658\,
            in2 => \N__9686\,
            in3 => \N__13592\,
            lcout => OPEN,
            ltout => \resetGen.reset_count_2_i_0_a3_5Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_i_0_a3_4_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8478\,
            in1 => \N__8472\,
            in2 => \N__8502\,
            in3 => \N__9969\,
            lcout => \resetGen.N_133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_5_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9682\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13524\,
            ce => \N__13570\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_7_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8466\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13524\,
            ce => \N__13570\,
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_i_0_a3_6_4_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13615\,
            in1 => \N__10009\,
            in2 => \N__9614\,
            in3 => \N__10063\,
            lcout => \resetGen.reset_count_2_i_0_a3_6Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_i_0_a3_4_4_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__10114\,
            in1 => \N__9713\,
            in2 => \_gnd_net_\,
            in3 => \N__9634\,
            lcout => \resetGen.reset_count_2_i_0_a3_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_1_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8451\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNI8RI7_0_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__10113\,
            in1 => \N__10072\,
            in2 => \N__10030\,
            in3 => \N__9970\,
            lcout => \buart.Z_rx.N_129\,
            ltout => \buart.Z_rx.N_129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_RNIVHME_0_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8465\,
            in2 => \N__8454\,
            in3 => \N__8450\,
            lcout => \buart.Z_rx.startbit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.Lab3U00.q_esr_ctle_7_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9945\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15917\,
            lcout => \Lab_UT.Lab3U00.bu_rx_data_rdy_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNIGM5F_0_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9944\,
            in2 => \_gnd_net_\,
            in3 => \N__9911\,
            lcout => \buart.Z_rx.N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec1.segmentUQ_0_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__14198\,
            in1 => \N__17335\,
            in2 => \N__14120\,
            in3 => \N__15646\,
            lcout => \L3_segment2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dicfsm.cState_RNO_3_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__8858\,
            in1 => \N__10364\,
            in2 => \N__8820\,
            in3 => \N__10316\,
            lcout => \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dek.det_N_0_a3_1_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8857\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8816\,
            lcout => \Lab_UT.dictrluu0.N_103_1\,
            ltout => \Lab_UT.dictrluu0.N_103_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dicfsm.cState_RNO_1_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10365\,
            in1 => \N__10312\,
            in2 => \N__8784\,
            in3 => \N__8781\,
            lcout => \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec3.g0_0_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000100000010"
        )
    port map (
            in0 => \N__15187\,
            in1 => \N__17061\,
            in2 => \N__15102\,
            in3 => \N__17450\,
            lcout => \N_52_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_3_1_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10182\,
            in1 => \N__8743\,
            in2 => \_gnd_net_\,
            in3 => \N__8575\,
            lcout => \uu2.un1_w_user_lf_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_44_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8744\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10183\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_26_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_31_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000001000"
        )
    port map (
            in0 => \N__12427\,
            in1 => \N__8667\,
            in2 => \N__8580\,
            in3 => \N__8576\,
            lcout => \uu2.mem0.G_14_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.Lab3U00.q_esr_1_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13626\,
            lcout => \Lab_UT_rx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13501\,
            ce => \N__9082\,
            sr => \N__15876\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12428\,
            in1 => \N__9048\,
            in2 => \_gnd_net_\,
            in3 => \N__11703\,
            lcout => \uu2.mem0.w_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI80631_4_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13995\,
            in2 => \_gnd_net_\,
            in3 => \N__13002\,
            lcout => \uu2.N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12840\,
            in1 => \N__8994\,
            in2 => \_gnd_net_\,
            in3 => \N__12429\,
            lcout => \uu2.mem0.w_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec1.g0_i_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011111011"
        )
    port map (
            in0 => \N__17342\,
            in1 => \N__14199\,
            in2 => \N__14121\,
            in3 => \N__15653\,
            lcout => \L3_segment2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_32_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8917\,
            in2 => \_gnd_net_\,
            in3 => \N__16183\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_19_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111110"
        )
    port map (
            in0 => \N__9228\,
            in1 => \N__8949\,
            in2 => \N__8943\,
            in3 => \N__12471\,
            lcout => \uu2.mem0.G_14_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI6NLE_7_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13847\,
            in2 => \_gnd_net_\,
            in3 => \N__14246\,
            lcout => OPEN,
            ltout => \uu2.N_329_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIV60G2_2_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10377\,
            in1 => \N__11698\,
            in2 => \N__8934\,
            in3 => \N__14988\,
            lcout => \uu2.Z_decfrac105_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_57_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__13791\,
            in1 => \N__9153\,
            in2 => \_gnd_net_\,
            in3 => \N__9144\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_2159_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_50_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14340\,
            in2 => \N__9138\,
            in3 => \N__13665\,
            lcout => \uu2.mem0.N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_20_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000001000"
        )
    port map (
            in0 => \N__11715\,
            in1 => \N__9243\,
            in2 => \N__9195\,
            in3 => \N__10414\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI0OT22_4_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__9180\,
            in1 => \N__9129\,
            in2 => \_gnd_net_\,
            in3 => \N__12657\,
            lcout => \uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4\,
            ltout => \uu2.w_addr_displaying_fast_RNI0OT22Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_41_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9186\,
            in2 => \N__9120\,
            in3 => \N__14425\,
            lcout => \uu2.mem0.un1_segment3_m2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_28_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__11597\,
            in1 => \N__10547\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_16_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011101111"
        )
    port map (
            in0 => \N__10500\,
            in1 => \N__9117\,
            in2 => \N__9111\,
            in3 => \N__10413\,
            lcout => \uu2.mem0.bitmap_pmux_1_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_38_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000001"
        )
    port map (
            in0 => \N__11596\,
            in1 => \N__12732\,
            in2 => \N__12645\,
            in3 => \N__9102\,
            lcout => \uu2.mem0.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_46_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9267\,
            in1 => \N__14426\,
            in2 => \_gnd_net_\,
            in3 => \N__10526\,
            lcout => \uu2.mem0.un1_segment3_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_27_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110111"
        )
    port map (
            in0 => \N__10548\,
            in1 => \N__11598\,
            in2 => \N__10418\,
            in3 => \N__10386\,
            lcout => \uu2.mem0.un1_segment3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_34_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__11589\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10546\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIHKAF2_0_8_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15366\,
            in1 => \N__12565\,
            in2 => \N__9279\,
            in3 => \N__12819\,
            lcout => \uu2.Z_decfrac106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_47_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111010"
        )
    port map (
            in0 => \N__12644\,
            in1 => \N__14400\,
            in2 => \N__12728\,
            in3 => \N__11588\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_35_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9204\,
            in2 => \N__9198\,
            in3 => \N__9171\,
            lcout => \uu2.mem0.un1_segment3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_55_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101111001"
        )
    port map (
            in0 => \N__16682\,
            in1 => \N__16966\,
            in2 => \N__16784\,
            in3 => \N__16875\,
            lcout => \uu2.mem0.N_2160_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec3.segmentUQ_i_0_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100100010000"
        )
    port map (
            in0 => \N__17064\,
            in1 => \N__15095\,
            in2 => \N__15189\,
            in3 => \N__17449\,
            lcout => \N_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_48_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__12643\,
            in1 => \N__14399\,
            in2 => \N__12727\,
            in3 => \N__11587\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_7_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11234\,
            in1 => \N__9165\,
            in2 => \_gnd_net_\,
            in3 => \N__9384\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13487\,
            ce => \N__9560\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_8_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9390\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11233\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13487\,
            ce => \N__9560\,
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__12470\,
            in1 => \_gnd_net_\,
            in2 => \N__9378\,
            in3 => \N__13782\,
            lcout => \uu2.mem0.w_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12469\,
            in1 => \N__9327\,
            in2 => \_gnd_net_\,
            in3 => \N__12293\,
            lcout => \uu2.mem0.w_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI362A1_3_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__15365\,
            in1 => \N__12796\,
            in2 => \_gnd_net_\,
            in3 => \N__14463\,
            lcout => \uu2.w_addr_displaying_RNI362A1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI50L01_0_2_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__11694\,
            in1 => \N__16193\,
            in2 => \_gnd_net_\,
            in3 => \N__14975\,
            lcout => \uu2.Z_decfrac106_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_56_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__16971\,
            in1 => \N__16874\,
            in2 => \N__16788\,
            in3 => \N__16683\,
            lcout => \uu2.mem0.N_2160_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9430\,
            in2 => \N__9411\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_1_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9462\,
            in3 => \N__9255\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__13540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10672\,
            in1 => \N__9449\,
            in2 => \_gnd_net_\,
            in3 => \N__9252\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__13540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9489\,
            in3 => \N__9510\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__13540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__10673\,
            in1 => \_gnd_net_\,
            in2 => \N__9501\,
            in3 => \N__9507\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__13540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__9476\,
            in1 => \N__10671\,
            in2 => \_gnd_net_\,
            in3 => \N__9504\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13540\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9497\,
            in1 => \N__9485\,
            in2 => \N__9477\,
            in3 => \N__9458\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__9406\,
            in1 => \N__9429\,
            in2 => \N__9450\,
            in3 => \N__9438\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_0_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100000010"
        )
    port map (
            in0 => \N__10670\,
            in1 => \N__10812\,
            in2 => \N__11189\,
            in3 => \N__10700\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9431\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__9432\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9410\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13532\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__10715\,
            in1 => \N__10811\,
            in2 => \_gnd_net_\,
            in3 => \N__10669\,
            lcout => \buart.Z_tx.un1_bitcount_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9527\,
            in2 => \N__9762\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9732\,
            in2 => \_gnd_net_\,
            in3 => \N__9591\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9889\,
            in1 => \N__9540\,
            in2 => \_gnd_net_\,
            in3 => \N__9588\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__13527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9791\,
            in2 => \_gnd_net_\,
            in3 => \N__9585\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__9777\,
            in1 => \N__9934\,
            in2 => \N__9896\,
            in3 => \N__9582\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__9792\,
            in1 => \N__9935\,
            in2 => \N__9579\,
            in3 => \N__9879\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13527\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIV5CT5_3_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10674\,
            in1 => \N__11922\,
            in2 => \_gnd_net_\,
            in3 => \N__10815\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9760\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9871\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9870\,
            in1 => \N__9526\,
            in2 => \_gnd_net_\,
            in3 => \N__9761\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9539\,
            in1 => \N__9730\,
            in2 => \N__9528\,
            in3 => \N__9790\,
            lcout => OPEN,
            ltout => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9776\,
            in2 => \N__9765\,
            in3 => \N__9759\,
            lcout => \buart.Z_rx.ser_clk\,
            ltout => \buart.Z_rx.ser_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__9741\,
            in1 => \N__9731\,
            in2 => \N__9735\,
            in3 => \N__9872\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000001"
        )
    port map (
            in0 => \N__10838\,
            in1 => \N__10881\,
            in2 => \N__10956\,
            in3 => \N__10962\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13521\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_6_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9709\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13513\,
            ce => \N__13577\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9659\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13513\,
            ce => \N__13577\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_2_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9610\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13513\,
            ce => \N__13577\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_3_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9635\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13513\,
            ce => \N__13577\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dek.det_N_0_o2_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__10195\,
            in1 => \N__10159\,
            in2 => \N__10128\,
            in3 => \N__10226\,
            lcout => \Lab_UT.dictrluu0.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dicfsm.cState_RNO_0_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10227\,
            in1 => \N__10196\,
            in2 => \N__10164\,
            in3 => \N__10127\,
            lcout => \Lab_UT.dictrluu0.dicfsm.nState_i_m3_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.Lab3U01.q_0_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10116\,
            in1 => \N__10074\,
            in2 => \N__10032\,
            in3 => \N__9972\,
            lcout => \Lab_UT.rx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13505\,
            ce => 'H',
            sr => \N__15882\
        );

    \buart.Z_rx.bitcount_e_0_RNI8RI7_0_0_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10115\,
            in1 => \N__10073\,
            in2 => \N__10031\,
            in3 => \N__9971\,
            lcout => bu_rx_data_rdy,
            ltout => \bu_rx_data_rdy_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_e_0_RNII0231_0_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__9936\,
            in1 => \N__9912\,
            in2 => \N__9900\,
            in3 => \N__9845\,
            lcout => \buart.Z_rx.bitcount_e_0_RNII0231Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec3.segmentUQ_0_6_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111101110"
        )
    port map (
            in0 => \N__15131\,
            in1 => \N__17003\,
            in2 => \N__17421\,
            in3 => \N__15047\,
            lcout => OPEN,
            ltout => \Lab_UT_dec3_segmentUQ_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment4_1_am_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__15049\,
            in1 => \N__9801\,
            in2 => \N__9804\,
            in3 => \N__15133\,
            lcout => \uu2.un1_segment4_1_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpmtens.q_RNIRE5_1_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17002\,
            in2 => \_gnd_net_\,
            in3 => \N__17393\,
            lcout => \N_71\,
            ltout => \N_71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpmtens.q_2_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001100"
        )
    port map (
            in0 => \N__10491\,
            in1 => \N__13152\,
            in2 => \N__9795\,
            in3 => \N__15134\,
            lcout => \Lab_UT_di_Mtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13500\,
            ce => 'H',
            sr => \N__15880\
        );

    \Lab_UT.dec3.segmentUQ_1_1_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010111110111"
        )
    port map (
            in0 => \N__15130\,
            in1 => \N__17005\,
            in2 => \N__17422\,
            in3 => \N__15046\,
            lcout => OPEN,
            ltout => \Lab_UT_dec3_segmentUQ_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment4_0_bm_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__15048\,
            in1 => \N__17400\,
            in2 => \N__10380\,
            in3 => \N__11406\,
            lcout => \uu2.un1_segment4_0_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpmtens.q_RNITG5_1_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__15132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17004\,
            lcout => \N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIAPHB1_0_5_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13771\,
            in1 => \N__12213\,
            in2 => \N__12315\,
            in3 => \N__12838\,
            lcout => \uu2.Z_decfrac105_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNID8KP2_2_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__12839\,
            in1 => \N__11699\,
            in2 => \N__12156\,
            in3 => \N__10455\,
            lcout => \uu2.g0_i_o4_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_1_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__17143\,
            in1 => \N__17080\,
            in2 => \_gnd_net_\,
            in3 => \N__10275\,
            lcout => \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dek.det_N_0_a3_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10262\,
            in1 => \N__10371\,
            in2 => \N__10320\,
            in3 => \N__10281\,
            lcout => \Lab_UT.dicSelectLEDdisp\,
            ltout => \Lab_UT.dicSelectLEDdisp_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_0_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__17079\,
            in1 => \_gnd_net_\,
            in2 => \N__10266\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.didpuu0.ledDisp00.selLedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dicfsm.cState_RNO_2_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__10263\,
            in1 => \N__10251\,
            in2 => \_gnd_net_\,
            in3 => \N__16569\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrluu0.dicfsm.N_102_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrluu0.dicfsm.cState_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__10245\,
            in1 => \N__10236\,
            in2 => \N__10230\,
            in3 => \N__15921\,
            lcout => \Lab_UT_dicRun\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIAGS21_4_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110101110"
        )
    port map (
            in0 => \N__13775\,
            in1 => \N__14462\,
            in2 => \N__14766\,
            in3 => \N__13996\,
            lcout => \uu2.un1_segment3_m4_s_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIU2OL2_5_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__13014\,
            in1 => \N__14510\,
            in2 => \N__11451\,
            in3 => \N__10454\,
            lcout => OPEN,
            ltout => \uu2.N_49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI9HV1J_5_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010111"
        )
    port map (
            in0 => \N__14472\,
            in1 => \N__12597\,
            in2 => \N__10443\,
            in3 => \N__10395\,
            lcout => \uu2.un1_segment3_m4_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIAH4P4_4_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__10440\,
            in1 => \N__11619\,
            in2 => \_gnd_net_\,
            in3 => \N__11466\,
            lcout => OPEN,
            ltout => \uu2.g0_i_o4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNINK1T81_2_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110010"
        )
    port map (
            in0 => \N__10434\,
            in1 => \N__10428\,
            in2 => \N__10422\,
            in3 => \N__11478\,
            lcout => \uu2.un1_segment3_m4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep1_RNIMMRIA_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12666\,
            in1 => \N__10464\,
            in2 => \_gnd_net_\,
            in3 => \N__11364\,
            lcout => \uu2.w_addr_displaying_4_rep1_RNIMMRIAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_53_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110111010"
        )
    port map (
            in0 => \N__12631\,
            in1 => \N__14398\,
            in2 => \N__11607\,
            in3 => \N__12731\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_53_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_40_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10515\,
            in2 => \N__10389\,
            in3 => \N__11508\,
            lcout => \uu2.mem0.un1_segment3_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_6_rep1_RNI9Q3H_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__14827\,
            in1 => \N__15457\,
            in2 => \_gnd_net_\,
            in3 => \N__16422\,
            lcout => \uu2.un1_segment4_sn_N_58_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_52_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15747\,
            in1 => \N__14427\,
            in2 => \_gnd_net_\,
            in3 => \N__10527\,
            lcout => \uu2.mem0.un1_segment3_m2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_42_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110111010"
        )
    port map (
            in0 => \N__12630\,
            in1 => \N__14397\,
            in2 => \N__11606\,
            in3 => \N__12730\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_30_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__10509\,
            in1 => \_gnd_net_\,
            in2 => \N__10503\,
            in3 => \N__11544\,
            lcout => \uu2.mem0.un1_segment3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec0.un137_segmentUQ_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14750\,
            in1 => \N__17246\,
            in2 => \N__14671\,
            in3 => \N__15729\,
            lcout => \Lab_UT_dec0_un137_segmentUQ\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment4_5_am_1_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100101010"
        )
    port map (
            in0 => \N__15730\,
            in1 => \N__14651\,
            in2 => \N__17255\,
            in3 => \N__14751\,
            lcout => \uu2.un1_segment4_5_amZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpmtens.q_RNO_0_2_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000100"
        )
    port map (
            in0 => \N__17448\,
            in1 => \N__15167\,
            in2 => \N__17063\,
            in3 => \N__15073\,
            lcout => \Lab_UT.didpuu0.didpmtens.q_5_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment4_1_bm_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010111101"
        )
    port map (
            in0 => \N__15166\,
            in1 => \N__17054\,
            in2 => \N__15088\,
            in3 => \N__17447\,
            lcout => OPEN,
            ltout => \uu2.un1_segment4_1_bmZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIPN54_8_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10479\,
            in2 => \N__10470\,
            in3 => \N__15248\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_fast_RNIPN54Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI9TKJ4_2_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13972\,
            in2 => \N__10467\,
            in3 => \N__10581\,
            lcout => \uu2.N_292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIV5694_2_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000010001"
        )
    port map (
            in0 => \N__10590\,
            in1 => \N__12868\,
            in2 => \N__10626\,
            in3 => \N__12954\,
            lcout => \uu2.w_addr_displaying_fast_RNIV5694Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIHV86_5_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__14568\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14511\,
            lcout => \uu2.N_290_0_i_0\,
            ltout => \uu2.N_290_0_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI1BU61_7_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__12795\,
            in1 => \N__13762\,
            in2 => \N__10575\,
            in3 => \N__16278\,
            lcout => OPEN,
            ltout => \uu2.un1_w_addr_displaying_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI90195_7_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__16279\,
            in1 => \N__10572\,
            in2 => \N__10566\,
            in3 => \N__16482\,
            lcout => \uu2.un1_w_addr_displaying_inv_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_51_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13770\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12812\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_39_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__12224\,
            in1 => \N__12291\,
            in2 => \N__10563\,
            in3 => \N__11595\,
            lcout => \uu2.mem0.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIAPHB1_5_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111101111111"
        )
    port map (
            in0 => \N__13769\,
            in1 => \N__12223\,
            in2 => \N__12305\,
            in3 => \N__12811\,
            lcout => \uu2.un1_segment3_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_5_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__12292\,
            in1 => \_gnd_net_\,
            in2 => \N__13916\,
            in3 => \N__16103\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_5C_net\,
            ce => 'H',
            sr => \N__15854\
        );

    \uu2.w_addr_displaying_3_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__12813\,
            in1 => \N__15492\,
            in2 => \_gnd_net_\,
            in3 => \N__16102\,
            lcout => \uu2.w_addr_displayingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_5C_net\,
            ce => 'H',
            sr => \N__15854\
        );

    \uu2.w_addr_displaying_0_rep1_RNIUUGB1_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000100"
        )
    port map (
            in0 => \N__11460\,
            in1 => \N__12810\,
            in2 => \N__13780\,
            in3 => \N__14312\,
            lcout => \uu2.un1_segment4_sn_N_38_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment4_2_bm_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110101010111"
        )
    port map (
            in0 => \N__14744\,
            in1 => \N__17248\,
            in2 => \N__14674\,
            in3 => \N__15732\,
            lcout => \uu2.un1_segment4_2_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.g1_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101111100"
        )
    port map (
            in0 => \N__15733\,
            in1 => \N__14745\,
            in2 => \N__17256\,
            in3 => \N__14664\,
            lcout => \uu2.gZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment4_5_bm_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__14743\,
            in1 => \N__17247\,
            in2 => \N__14673\,
            in3 => \N__15731\,
            lcout => \uu2.un1_segment4_5_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_RNO_0_3_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111011101"
        )
    port map (
            in0 => \N__15734\,
            in1 => \N__14747\,
            in2 => \_gnd_net_\,
            in3 => \N__17253\,
            lcout => \Lab_UT.didpuu0.didpsones.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_RNI0GG11_3_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__14746\,
            in1 => \_gnd_net_\,
            in2 => \N__14675\,
            in3 => \N__17252\,
            lcout => \Lab_UT.didpuu0.didpsones.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMU_0_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17093\,
            in1 => \N__14191\,
            in2 => \_gnd_net_\,
            in3 => \N__14748\,
            lcout => OPEN,
            ltout => \Lab_UT.didpuu0.ledDisp00.selLed_RNIGTMUZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNIEH0Q1_1_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__17150\,
            in1 => \_gnd_net_\,
            in2 => \N__10614\,
            in3 => \N__10596\,
            lcout => led_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJ_0_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17094\,
            in1 => \N__16970\,
            in2 => \_gnd_net_\,
            in3 => \N__15188\,
            lcout => \Lab_UT.didpuu0.ledDisp00.selLed_RNIR2SJZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.un1_bitcount_cry_0_c_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10632\,
            in2 => \N__10701\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_2_0_\,
            carryout => \buart.Z_tx.un1_bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_1_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__11164\,
            in1 => \N__10755\,
            in2 => \N__10731\,
            in3 => \N__10776\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \buart.Z_tx.un1_bitcount_cry_0\,
            carryout => \buart.Z_tx.un1_bitcount_cry_1\,
            clk => \N__13543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_2_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__11165\,
            in1 => \N__10761\,
            in2 => \N__10749\,
            in3 => \N__10773\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.un1_bitcount_cry_1\,
            carryout => \buart.Z_tx.un1_bitcount_cry_2\,
            clk => \N__13543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_3_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111101110"
        )
    port map (
            in0 => \N__10770\,
            in1 => \N__11166\,
            in2 => \_gnd_net_\,
            in3 => \N__10764\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13543\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIM5O32_2_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__10668\,
            in1 => \_gnd_net_\,
            in2 => \N__10813\,
            in3 => \N__10748\,
            lcout => \buart.Z_tx.bitcount_RNIM5O32Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIL4O32_1_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \N__10730\,
            in1 => \N__10801\,
            in2 => \_gnd_net_\,
            in3 => \N__10667\,
            lcout => \buart.Z_tx.bitcount_RNIL4O32Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIQOQA1_3_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10744\,
            in1 => \N__10726\,
            in2 => \N__10716\,
            in3 => \N__10695\,
            lcout => \buart__tx_uart_busy_0\,
            ltout => \buart__tx_uart_busy_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.un1_bitcount_cry_0_c_RNO_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \N__10696\,
            in1 => \_gnd_net_\,
            in2 => \N__10677\,
            in3 => \N__10666\,
            lcout => \buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_8_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__12101\,
            in1 => \N__12009\,
            in2 => \_gnd_net_\,
            in3 => \N__12077\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13537\,
            ce => 'H',
            sr => \N__15890\
        );

    \resetGen.reset_count_RNITEEC1_2_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__10905\,
            in1 => \N__10891\,
            in2 => \_gnd_net_\,
            in3 => \N__10823\,
            lcout => \resetGen.N_117\,
            ltout => \resetGen.N_117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001110"
        )
    port map (
            in0 => \N__10955\,
            in1 => \N__10880\,
            in2 => \N__10941\,
            in3 => \N__10851\,
            lcout => \resetGen.reset_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__10849\,
            in1 => \N__10878\,
            in2 => \N__10911\,
            in3 => \N__10893\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__10877\,
            in1 => \N__10907\,
            in2 => \_gnd_net_\,
            in3 => \N__10848\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10876\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNO_0_2_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__10906\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10892\,
            lcout => OPEN,
            ltout => \resetGen.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101001"
        )
    port map (
            in0 => \N__10824\,
            in1 => \N__10879\,
            in2 => \N__10854\,
            in3 => \N__10850\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13530\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_10__un382_ci_8_1_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12131\,
            in1 => \N__11952\,
            in2 => \N__12054\,
            in3 => \N__11977\,
            lcout => \uu2.vbuf_count.un382_ci_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_7__un349_ci_0_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11978\,
            in1 => \N__12052\,
            in2 => \_gnd_net_\,
            in3 => \N__11953\,
            lcout => \uu2.un349_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIQF5F5_4_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10814\,
            in2 => \_gnd_net_\,
            in3 => \N__11913\,
            lcout => vbuf_tx_data_rdy,
            ltout => \vbuf_tx_data_rdy_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIU80H5_4_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11355\,
            in3 => \N__15920\,
            lcout => \uu2.vbuf_tx_data_rdy_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_4_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__12053\,
            in1 => \N__12017\,
            in2 => \_gnd_net_\,
            in3 => \N__11914\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13525\,
            ce => 'H',
            sr => \N__15886\
        );

    \uu2.r_addr_1_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11279\,
            in1 => \N__11304\,
            in2 => \_gnd_net_\,
            in3 => \N__11162\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13525\,
            ce => 'H',
            sr => \N__15886\
        );

    \uu2.r_addr_2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11305\,
            in1 => \N__11272\,
            in2 => \N__11103\,
            in3 => \N__11163\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13518\,
            ce => 'H',
            sr => \N__15884\
        );

    \Lab_UT.didpuu0.didpmtens.q_0_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__13215\,
            in1 => \N__13183\,
            in2 => \_gnd_net_\,
            in3 => \N__17420\,
            lcout => \Lab_UT_di_Mtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13511\,
            ce => 'H',
            sr => \N__15883\
        );

    \uu2.un1_segment4_2_am_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12240\,
            in2 => \_gnd_net_\,
            in3 => \N__12872\,
            lcout => \uu2.un1_segment4_2_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.sec_clk_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11076\,
            in2 => \_gnd_net_\,
            in3 => \N__16537\,
            lcout => \Lab_UT_l_oneSecPluse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13511\,
            ce => 'H',
            sr => \N__15883\
        );

    \Lab_UT.secuu0.delay_line_1_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10995\,
            lcout => \Lab_UT.secuu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13511\,
            ce => 'H',
            sr => \N__15883\
        );

    \Lab_UT.didpuu0.didpmtens.q_1_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011001001100"
        )
    port map (
            in0 => \N__13151\,
            in1 => \N__17045\,
            in2 => \N__11418\,
            in3 => \N__17419\,
            lcout => \Lab_UT_di_Mtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13502\,
            ce => 'H',
            sr => \N__15879\
        );

    \Lab_UT.didpuu0.didpmtens.q_RNO_0_1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17417\,
            in1 => \N__15051\,
            in2 => \_gnd_net_\,
            in3 => \N__15137\,
            lcout => \Lab_UT.didpuu0.didpmtens.N_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec3.segmentUQ_0_o2_5_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__15135\,
            in1 => \N__17043\,
            in2 => \_gnd_net_\,
            in3 => \N__17415\,
            lcout => OPEN,
            ltout => \N_84_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment4_0_am_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001110011"
        )
    port map (
            in0 => \N__17416\,
            in1 => \N__15050\,
            in2 => \N__11409\,
            in3 => \N__11405\,
            lcout => OPEN,
            ltout => \uu2.un1_segment4_0_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIK7I7_2_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000111"
        )
    port map (
            in0 => \N__11394\,
            in1 => \N__12962\,
            in2 => \N__11388\,
            in3 => \N__12988\,
            lcout => OPEN,
            ltout => \uu2.un1_segment4_8_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep1_RNI6JSF4_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__11385\,
            in1 => \N__14822\,
            in2 => \N__11373\,
            in3 => \N__11370\,
            lcout => \uu2.N_286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec3.un75_segmentUQ_i_i_o2_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__15136\,
            in1 => \N__17044\,
            in2 => \_gnd_net_\,
            in3 => \N__17418\,
            lcout => OPEN,
            ltout => \Lab_UT.N_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpmtens.q_3_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__13184\,
            in1 => \N__13214\,
            in2 => \N__11358\,
            in3 => \N__15052\,
            lcout => \Lab_UT_di_Mtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13502\,
            ce => 'H',
            sr => \N__15879\
        );

    \uu2.w_addr_displaying_fast_RNIK9D9_2_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12952\,
            in1 => \N__14554\,
            in2 => \_gnd_net_\,
            in3 => \N__13060\,
            lcout => \uu2.un1_segment4_sn_N_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNILAD9_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__14555\,
            in1 => \N__12953\,
            in2 => \_gnd_net_\,
            in3 => \N__12989\,
            lcout => OPEN,
            ltout => \uu2.g0_i_o4_0_a8_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_5_rep1_RNIVO2E1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__12924\,
            in1 => \N__13851\,
            in2 => \N__11469\,
            in3 => \N__16473\,
            lcout => \uu2.w_addr_displaying_5_rep1_RNIVO2EZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_4_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__15292\,
            in1 => \_gnd_net_\,
            in2 => \N__16092\,
            in3 => \N__12990\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_4C_net\,
            ce => 'H',
            sr => \N__15850\
        );

    \uu2.w_addr_displaying_fast_6_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16049\,
            in2 => \N__12585\,
            in3 => \N__14556\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_4C_net\,
            ce => 'H',
            sr => \N__15850\
        );

    \uu2.w_addr_displaying_8_rep1_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__13852\,
            in1 => \N__16059\,
            in2 => \N__15306\,
            in3 => \N__15369\,
            lcout => \uu2.w_addr_displaying_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_4C_net\,
            ce => 'H',
            sr => \N__15850\
        );

    \uu2.w_addr_displaying_8_rep1_RNIN6OC_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__13826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14887\,
            lcout => \uu2.N_315_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_7_rep1_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__14888\,
            in1 => \N__16058\,
            in2 => \N__13913\,
            in3 => \N__14013\,
            lcout => \uu2.w_addr_displaying_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_4C_net\,
            ce => 'H',
            sr => \N__15850\
        );

    \uu2.w_addr_displaying_2_rep1_RNIQ3R01_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__15458\,
            in1 => \N__14307\,
            in2 => \N__15552\,
            in3 => \N__16365\,
            lcout => \uu2.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep2_RNI5R4M_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010011001"
        )
    port map (
            in0 => \N__14308\,
            in1 => \N__11685\,
            in2 => \_gnd_net_\,
            in3 => \N__15551\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_1_1_3_tz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIDUPM1_2_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110011111"
        )
    port map (
            in0 => \N__11686\,
            in1 => \N__12834\,
            in2 => \N__11442\,
            in3 => \N__14999\,
            lcout => \uu2.bitmap_pmux_1_1_3_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI50L01_2_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11687\,
            in1 => \N__16184\,
            in2 => \_gnd_net_\,
            in3 => \N__15000\,
            lcout => \uu2.N_111\,
            ltout => \uu2.N_111_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.counter_gen_label_5__un436_ci_0_a2_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__12835\,
            in1 => \_gnd_net_\,
            in2 => \N__11523\,
            in3 => \N__13757\,
            lcout => \uu2.un436_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__13758\,
            in1 => \N__15291\,
            in2 => \_gnd_net_\,
            in3 => \N__16083\,
            lcout => \uu2.w_addr_displayingZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__15852\
        );

    \uu2.w_addr_displaying_fast_2_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__16082\,
            in1 => \N__15001\,
            in2 => \N__16199\,
            in3 => \N__12961\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__15852\
        );

    \uu2.w_addr_displaying_5_rep1_RNI50LS_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16421\,
            in1 => \N__15459\,
            in2 => \N__14902\,
            in3 => \N__16472\,
            lcout => OPEN,
            ltout => \uu2.un1_segment4_sn_N_36_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_5_rep1_RNIMG8P2_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__16547\,
            in1 => \N__16570\,
            in2 => \N__11520\,
            in3 => \N__11517\,
            lcout => \uu2.N_2150_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_54_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010000"
        )
    port map (
            in0 => \N__14386\,
            in1 => \N__12618\,
            in2 => \N__11599\,
            in3 => \N__12715\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIKR5D1_6_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111111111"
        )
    port map (
            in0 => \N__12222\,
            in1 => \N__11502\,
            in2 => \N__12575\,
            in3 => \N__13983\,
            lcout => OPEN,
            ltout => \uu2.g2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_rep1_RNIN998E_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__11496\,
            in1 => \N__11490\,
            in2 => \N__11481\,
            in3 => \N__13089\,
            lcout => \uu2.N_299_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_43_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010000"
        )
    port map (
            in0 => \N__12617\,
            in1 => \N__14385\,
            in2 => \N__12729\,
            in3 => \N__11586\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIUCHB1_3_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15480\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12837\,
            lcout => \uu2.un15_w_data_displaying_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec2.segmentUQ_2_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111111011"
        )
    port map (
            in0 => \N__16670\,
            in1 => \N__16859\,
            in2 => \N__16965\,
            in3 => \N__16721\,
            lcout => \L3_segment3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpmones.q_esr_3_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110100011110000"
        )
    port map (
            in0 => \N__16863\,
            in1 => \N__16953\,
            in2 => \N__16743\,
            in3 => \N__16674\,
            lcout => \Lab_UT_di_Mones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13488\,
            ce => \N__11865\,
            sr => \N__15887\
        );

    \uu2.segment3_m_1_6_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101111100"
        )
    port map (
            in0 => \N__16672\,
            in1 => \N__16861\,
            in2 => \N__16964\,
            in3 => \N__16720\,
            lcout => OPEN,
            ltout => \uu2.segment3_m_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_7_rep1_RNIA86H1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11538\,
            in3 => \N__14892\,
            lcout => OPEN,
            ltout => \uu2.segment3_m_2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIE28D2_4_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__13763\,
            in1 => \N__12794\,
            in2 => \N__11535\,
            in3 => \N__13973\,
            lcout => \uu2.segment3_m_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment4_4_bm_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011111011"
        )
    port map (
            in0 => \N__16860\,
            in1 => \N__16946\,
            in2 => \N__16742\,
            in3 => \N__16671\,
            lcout => \uu2.un1_segment4_4_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment4_4_am_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101110001"
        )
    port map (
            in0 => \N__16673\,
            in1 => \N__16862\,
            in2 => \N__16963\,
            in3 => \N__16716\,
            lcout => OPEN,
            ltout => \uu2.un1_segment4_4_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNICB763_0_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__15249\,
            in1 => \N__11532\,
            in2 => \N__11526\,
            in3 => \N__15944\,
            lcout => \uu2.un1_segment4_9_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_23_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__12571\,
            in1 => \N__11736\,
            in2 => \N__12483\,
            in3 => \N__16285\,
            lcout => \uu2.mem0.G_14_0_a6_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_36_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101111110111"
        )
    port map (
            in0 => \N__12799\,
            in1 => \N__11662\,
            in2 => \N__11730\,
            in3 => \N__14993\,
            lcout => \uu2.mem0.bitmap_pmux_1_1_2_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI83L01_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111010"
        )
    port map (
            in0 => \N__13765\,
            in1 => \_gnd_net_\,
            in2 => \N__11684\,
            in3 => \N__16175\,
            lcout => \uu2.bitmap_pmux_1_1_2_tz_1_0\,
            ltout => \uu2.bitmap_pmux_1_1_2_tz_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_45_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101111110111"
        )
    port map (
            in0 => \N__12798\,
            in1 => \N__11661\,
            in2 => \N__11721\,
            in3 => \N__14992\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_1_1_2_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_33_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__12570\,
            in1 => \_gnd_net_\,
            in2 => \N__11718\,
            in3 => \N__16284\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__16176\,
            in1 => \N__11663\,
            in2 => \N__16104\,
            in3 => \N__14994\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2C_net\,
            ce => 'H',
            sr => \N__15857\
        );

    \uu2.w_addr_displaying_RNI8NHB1_2_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110101"
        )
    port map (
            in0 => \N__13764\,
            in1 => \N__12797\,
            in2 => \N__11683\,
            in3 => \N__16283\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_RNI8NHB1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI18582_8_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001010111010"
        )
    port map (
            in0 => \N__13020\,
            in1 => \N__12569\,
            in2 => \N__11622\,
            in3 => \N__13997\,
            lcout => \uu2.w_addr_displaying_RNI18582Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec2.un152_segmentUQ_1_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16754\,
            in2 => \_gnd_net_\,
            in3 => \N__16939\,
            lcout => \Lab_UT.un152_segmentUQ_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI89GK1_2_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__11955\,
            in1 => \N__11841\,
            in2 => \N__12078\,
            in3 => \N__11821\,
            lcout => \uu2.un3_r_clk_en_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_2_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__11783\,
            in1 => \N__11825\,
            in2 => \N__11849\,
            in3 => \N__11921\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13544\,
            ce => 'H',
            sr => \N__15893\
        );

    \uu2.l_count_0_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11822\,
            in2 => \_gnd_net_\,
            in3 => \N__11919\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13544\,
            ce => 'H',
            sr => \N__15893\
        );

    \uu2.l_count_3_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11784\,
            in1 => \N__11848\,
            in2 => \N__11802\,
            in3 => \N__11826\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13544\,
            ce => 'H',
            sr => \N__15893\
        );

    \uu2.vbuf_count.counter_gen_label_4__un316_ci_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11823\,
            in1 => \N__11798\,
            in2 => \N__11850\,
            in3 => \N__11781\,
            lcout => \uu2.un316_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_1_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11782\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11824\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13544\,
            ce => 'H',
            sr => \N__15893\
        );

    \uu2.l_count_RNI89GK1_3_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__11975\,
            in1 => \N__11797\,
            in2 => \N__12132\,
            in3 => \N__11780\,
            lcout => \uu2.un3_r_clk_en_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI626E_10_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11879\,
            in2 => \_gnd_net_\,
            in3 => \N__12112\,
            lcout => OPEN,
            ltout => \uu2.un3_r_clk_en_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI0NA44_4_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12039\,
            in1 => \N__11763\,
            in2 => \N__11757\,
            in3 => \N__11754\,
            lcout => uu2_un3_r_clk_en_0,
            ltout => \uu2_un3_r_clk_en_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_5_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__11976\,
            in1 => \N__12008\,
            in2 => \N__12144\,
            in3 => \N__12040\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13538\,
            ce => 'H',
            sr => \N__15892\
        );

    \uu2.l_count_7_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__12006\,
            in1 => \N__12130\,
            in2 => \N__12141\,
            in3 => \N__11918\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13538\,
            ce => 'H',
            sr => \N__15892\
        );

    \uu2.l_count_9_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12076\,
            in1 => \N__12007\,
            in2 => \N__12102\,
            in3 => \N__12114\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13538\,
            ce => 'H',
            sr => \N__15892\
        );

    \uu2.vbuf_count.counter_gen_label_10__un382_ci_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12113\,
            in1 => \N__12097\,
            in2 => \N__12016\,
            in3 => \N__12075\,
            lcout => \uu2.un382_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_6_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__12048\,
            in1 => \N__11954\,
            in2 => \N__12021\,
            in3 => \N__11979\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13531\,
            ce => 'H',
            sr => \N__15889\
        );

    \uu2.l_count_10_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__11928\,
            in1 => \N__11880\,
            in2 => \_gnd_net_\,
            in3 => \N__11920\,
            lcout => \uu2.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13531\,
            ce => 'H',
            sr => \N__15889\
        );

    \Lab_UT.didpuu0.didpstens.q_RNIL3BL3_1_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__13177\,
            in1 => \N__17325\,
            in2 => \N__13244\,
            in3 => \N__15635\,
            lcout => \Lab_UT.didpuu0.countEnMones\,
            ltout => \Lab_UT.didpuu0.countEnMones_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpmones.q_esr_RNO_0_3_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11868\,
            in3 => \N__15918\,
            lcout => \Lab_UT.didpuu0.didpmones.countEnMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpstens.q_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011011001100"
        )
    port map (
            in0 => \N__13179\,
            in1 => \N__17326\,
            in2 => \N__13245\,
            in3 => \N__15637\,
            lcout => \Lab_UT_di_Stens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13519\,
            ce => 'H',
            sr => \N__15885\
        );

    \Lab_UT.didpuu0.didpstens.q_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15636\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13178\,
            lcout => \Lab_UT_di_Stens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13519\,
            ce => 'H',
            sr => \N__15885\
        );

    \Lab_UT.didpuu0.didpsones.q_RNIHCAV1_0_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15690\,
            in1 => \N__12917\,
            in2 => \_gnd_net_\,
            in3 => \N__13306\,
            lcout => \Lab_UT.didpuu0.countEnStens\,
            ltout => \Lab_UT.didpuu0.countEnStens_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpstens.q_esr_ctle_3_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12243\,
            in3 => \N__15919\,
            lcout => \Lab_UT.didpuu0.didpstens.countEnStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15691\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13307\,
            lcout => \Lab_UT_di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13519\,
            ce => 'H',
            sr => \N__15885\
        );

    \uu2.un1_segment4_2_am_1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100000100"
        )
    port map (
            in0 => \N__14734\,
            in1 => \N__17237\,
            in2 => \N__14672\,
            in3 => \N__15689\,
            lcout => \uu2.un1_segment4_2_amZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNO_0_6_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111011111010"
        )
    port map (
            in0 => \N__12338\,
            in1 => \N__12324\,
            in2 => \N__12225\,
            in3 => \N__13918\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_4_0_i_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_6_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12212\,
            in2 => \N__12234\,
            in3 => \N__16057\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_6C_net\,
            ce => 'H',
            sr => \N__15849\
        );

    \uu2.w_addr_displaying_RNIKFL01_6_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__12523\,
            in1 => \N__12181\,
            in2 => \_gnd_net_\,
            in3 => \N__13781\,
            lcout => \uu2.g0_i_o4_0_a8_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_8_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__12534\,
            in1 => \N__16056\,
            in2 => \N__15309\,
            in3 => \N__15346\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_6C_net\,
            ce => 'H',
            sr => \N__15849\
        );

    \uu2.w_addr_displaying_fast_RNO_0_6_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111011111010"
        )
    port map (
            in0 => \N__12337\,
            in1 => \N__12323\,
            in2 => \N__14573\,
            in3 => \N__13917\,
            lcout => \uu2.w_addr_displaying_4_0_i_fast_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIHKAF2_8_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15301\,
            in1 => \N__12524\,
            in2 => \_gnd_net_\,
            in3 => \N__15345\,
            lcout => \uu2.un15_w_data_displaying\,
            ltout => \uu2.un15_w_data_displaying_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIMF2HD_8_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12486\,
            in3 => \N__12426\,
            lcout => \uu2.un21_w_addr_displaying_i\,
            ltout => \uu2.un21_w_addr_displaying_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_7_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001101100"
        )
    port map (
            in0 => \N__13919\,
            in1 => \N__16251\,
            in2 => \N__12345\,
            in3 => \N__14012\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_6C_net\,
            ce => 'H',
            sr => \N__15849\
        );

    \uu2.w_addr_displaying_6_rep1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16045\,
            in1 => \N__12252\,
            in2 => \_gnd_net_\,
            in3 => \N__16414\,
            lcout => \uu2.w_addr_displaying_6_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_6_rep1C_net\,
            ce => 'H',
            sr => \N__15853\
        );

    \uu2.w_addr_displaying_6_rep1_RNO_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011111010"
        )
    port map (
            in0 => \N__16413\,
            in1 => \N__13914\,
            in2 => \N__12342\,
            in3 => \N__12316\,
            lcout => \uu2.w_addr_displaying_4_0_i_rep1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_5_rep1_RNI3HMT_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16409\,
            in1 => \N__16459\,
            in2 => \N__15456\,
            in3 => \N__15531\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_5_rep1_RNI3HMTZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_5_rep1_RNIMFM34_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13638\,
            in2 => \N__12246\,
            in3 => \N__14019\,
            lcout => \uu2.un1_segment3_m5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_5_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__13915\,
            in1 => \_gnd_net_\,
            in2 => \N__16091\,
            in3 => \N__14502\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_6_rep1C_net\,
            ce => 'H',
            sr => \N__15853\
        );

    \uu2.w_addr_displaying_fast_RNID5QH_5_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__14500\,
            in1 => \N__14557\,
            in2 => \_gnd_net_\,
            in3 => \N__13822\,
            lcout => \uu2.w_addr_displaying_fast_RNID5QHZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI6N2K_5_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__14558\,
            in1 => \N__14501\,
            in2 => \N__13843\,
            in3 => \N__15532\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_fast_RNI6N2KZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI76AF1_2_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__12681\,
            in1 => \_gnd_net_\,
            in2 => \N__12675\,
            in3 => \N__12672\,
            lcout => \uu2.un1_segment4_sn_N_39_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI2VHC_4_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__12986\,
            in1 => \N__13069\,
            in2 => \N__15247\,
            in3 => \N__14234\,
            lcout => \uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4\,
            ltout => \uu2.w_addr_displaying_fast_RNI2VHCZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNILB202_4_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__13756\,
            in1 => \N__13680\,
            in2 => \N__12648\,
            in3 => \N__14454\,
            lcout => \uu2.w_addr_displaying_RNILB202Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_rep1_RNIR94U_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010001010"
        )
    port map (
            in0 => \N__14453\,
            in1 => \N__15452\,
            in2 => \N__15546\,
            in3 => \N__16347\,
            lcout => \uu2.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep2_RNI75VM_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__13828\,
            in1 => \N__15426\,
            in2 => \N__14889\,
            in3 => \N__15533\,
            lcout => \uu2.w_addr_displaying_4_rep2_RNI75VMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_rep1_RNI4RA21_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15425\,
            in1 => \N__13827\,
            in2 => \N__16364\,
            in3 => \N__14866\,
            lcout => \uu2.un1_w_addr_displaying_inv_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_3_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13077\,
            in2 => \N__15490\,
            in3 => \N__16090\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_3C_net\,
            ce => 'H',
            sr => \N__15855\
        );

    \uu2.w_addr_displaying_fast_RNIN0TS_4_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__12985\,
            in1 => \N__14288\,
            in2 => \N__13082\,
            in3 => \N__16346\,
            lcout => \uu2.w_addr_displaying_fast_RNIN0TSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNILHHC_0_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__13070\,
            in1 => \N__12987\,
            in2 => \N__12963\,
            in3 => \N__15945\,
            lcout => \uu2.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpsones.q_1_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011001001100"
        )
    port map (
            in0 => \N__13321\,
            in1 => \N__17210\,
            in2 => \N__12918\,
            in3 => \N__15714\,
            lcout => \Lab_UT_di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13493\,
            ce => 'H',
            sr => \N__15888\
        );

    \Lab_UT.didpuu0.didpsones.q_2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__15715\,
            in1 => \N__13322\,
            in2 => \N__17238\,
            in3 => \N__14720\,
            lcout => \Lab_UT_di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13493\,
            ce => 'H',
            sr => \N__15888\
        );

    \Lab_UT.didpuu0.didpsones.q_3_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011000100"
        )
    port map (
            in0 => \N__13323\,
            in1 => \N__14619\,
            in2 => \N__12891\,
            in3 => \N__12873\,
            lcout => \Lab_UT_di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13493\,
            ce => 'H',
            sr => \N__15888\
        );

    \uu2.segment1_m_2_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__14719\,
            in1 => \N__17209\,
            in2 => \N__14637\,
            in3 => \N__15713\,
            lcout => OPEN,
            ltout => \uu2.segment1_m_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_7_rep1_RNIPUSD1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12846\,
            in3 => \N__14896\,
            lcout => OPEN,
            ltout => \uu2.segment1_m_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIBOM74_3_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__15367\,
            in1 => \N__13278\,
            in2 => \N__12843\,
            in3 => \N__12836\,
            lcout => OPEN,
            ltout => \uu2.un1_segment1_iv_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_rep1_RNI2NR6D_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__14319\,
            in1 => \N__12741\,
            in2 => \N__12735\,
            in3 => \N__16209\,
            lcout => \uu2.un1_segment1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpstens.q_esr_2_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011000100"
        )
    port map (
            in0 => \N__15640\,
            in1 => \N__14160\,
            in2 => \N__14090\,
            in3 => \N__17329\,
            lcout => \Lab_UT_di_Stens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13490\,
            ce => \N__13119\,
            sr => \N__15891\
        );

    \Lab_UT.didpuu0.didpstens.q_esr_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__15641\,
            in1 => \N__14161\,
            in2 => \N__14091\,
            in3 => \N__17330\,
            lcout => \Lab_UT_di_Stens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13490\,
            ce => \N__13119\,
            sr => \N__15891\
        );

    \uu2.un1_segment4_3_bm_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__14158\,
            in1 => \N__17327\,
            in2 => \N__14088\,
            in3 => \N__15638\,
            lcout => \uu2.un1_segment4_3_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment4_3_am_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110110111"
        )
    port map (
            in0 => \N__15639\,
            in1 => \N__14159\,
            in2 => \N__14089\,
            in3 => \N__17328\,
            lcout => OPEN,
            ltout => \uu2.un1_segment4_3_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_rep1_RNI8N8R6_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__14306\,
            in1 => \N__13107\,
            in2 => \N__13101\,
            in3 => \N__13098\,
            lcout => OPEN,
            ltout => \uu2.N_289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIFU9M8_8_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15561\,
            in1 => \_gnd_net_\,
            in2 => \N__13092\,
            in3 => \N__15195\,
            lcout => \uu2.w_addr_displaying_fast_RNIFU9M8Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIBHTT_3_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010110101001"
        )
    port map (
            in0 => \N__16363\,
            in1 => \N__13081\,
            in2 => \N__15002\,
            in3 => \N__14826\,
            lcout => \uu2.N_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep1_RNIAVDB_0_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__15450\,
            in1 => \_gnd_net_\,
            in2 => \N__14831\,
            in3 => \N__14906\,
            lcout => \uu2.w_addr_displaying_4_rep1_RNIAVDBZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIKFIE_6_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__15547\,
            in1 => \N__15451\,
            in2 => \N__14907\,
            in3 => \N__14574\,
            lcout => \uu2.w_addr_displaying_fast_RNIKFIEZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMU_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14071\,
            in1 => \N__14650\,
            in2 => \_gnd_net_\,
            in3 => \N__17111\,
            lcout => OPEN,
            ltout => \Lab_UT.didpuu0.ledDisp00.selLed_RNIIVMUZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNIRNGO1_1_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__13251\,
            in1 => \_gnd_net_\,
            in2 => \N__13266\,
            in3 => \N__17164\,
            lcout => led_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNI67CI_0_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17110\,
            in1 => \N__16741\,
            in2 => \_gnd_net_\,
            in3 => \N__15099\,
            lcout => \Lab_UT.didpuu0.ledDisp00.selLed_RNI67CIZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec1.un11_segmentUQ_1_0_a2_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14167\,
            in2 => \_gnd_net_\,
            in3 => \N__14070\,
            lcout => \Lab_UT.un11_segmentUQ_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpmones.q_esr_RNIF7VF1_3_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16930\,
            in1 => \N__16841\,
            in2 => \N__16782\,
            in3 => \N__16658\,
            lcout => OPEN,
            ltout => \Lab_UT.didpuu0.countEnMtens_0_a4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpstens.q_RNIJUV53_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__13229\,
            in1 => \N__17331\,
            in2 => \N__13218\,
            in3 => \N__15642\,
            lcout => \Lab_UT.didpuu0.countEnMtens_0_a4_1\,
            ltout => \Lab_UT.didpuu0.countEnMtens_0_a4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpstens.q_RNI4BA55_1_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13191\,
            in3 => \N__13188\,
            lcout => \Lab_UT.didpuu0.countEnMtens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpmones.q_2_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__16659\,
            in1 => \N__13656\,
            in2 => \N__16865\,
            in3 => \N__16931\,
            lcout => \Lab_UT_di_Mones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13485\,
            ce => 'H',
            sr => \N__15894\
        );

    \uu2.segment3_m_3_1_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110101010111"
        )
    port map (
            in0 => \N__16928\,
            in1 => \N__16840\,
            in2 => \N__16781\,
            in3 => \N__16657\,
            lcout => \uu2.segment3_m_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.didpmones.q_1_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010011110000"
        )
    port map (
            in0 => \N__13125\,
            in1 => \N__16668\,
            in2 => \N__16866\,
            in3 => \N__13655\,
            lcout => \Lab_UT_di_Mones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13485\,
            ce => 'H',
            sr => \N__15894\
        );

    \Lab_UT.didpuu0.didpmones.q_0_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13654\,
            in2 => \_gnd_net_\,
            in3 => \N__16660\,
            lcout => \Lab_UT_di_Mones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13485\,
            ce => 'H',
            sr => \N__15894\
        );

    \uu2.un1_segment3_m5_bm_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111010110101"
        )
    port map (
            in0 => \N__16656\,
            in1 => \N__16767\,
            in2 => \N__16864\,
            in3 => \N__16929\,
            lcout => \uu2.un1_segment3_m5_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13622\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13539\,
            ce => \N__13578\,
            sr => \_gnd_net_\
        );

    \Lab_UT.secuu0.sec_clkD_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16542\,
            lcout => \Lab_UT.sec_clkD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13526\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.clkSecStrb_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__16541\,
            in1 => \N__13334\,
            in2 => \_gnd_net_\,
            in3 => \N__16577\,
            lcout => \Lab_UT.didpuu0.clkSecStrbZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.segment2_m_2_5_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001011111011"
        )
    port map (
            in0 => \N__14187\,
            in1 => \N__17299\,
            in2 => \N__14110\,
            in3 => \N__15610\,
            lcout => \uu2.segment2_m_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec1.segmentUQ_4_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111010001"
        )
    port map (
            in0 => \N__15628\,
            in1 => \N__14190\,
            in2 => \N__14112\,
            in3 => \N__17317\,
            lcout => OPEN,
            ltout => \L3_segment2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep1_RNIBG883_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13293\,
            in2 => \N__13281\,
            in3 => \N__14791\,
            lcout => \uu2.un1_segment3_m0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.segment2_m_1_6_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110111100"
        )
    port map (
            in0 => \N__15627\,
            in1 => \N__14189\,
            in2 => \N__14111\,
            in3 => \N__17318\,
            lcout => \uu2.segment2_m_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_segment3_m5_am_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010111101"
        )
    port map (
            in0 => \N__14188\,
            in1 => \N__17316\,
            in2 => \N__14113\,
            in3 => \N__15626\,
            lcout => \uu2.un1_segment3_m5_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__14792\,
            in1 => \N__15305\,
            in2 => \_gnd_net_\,
            in3 => \N__16054\,
            lcout => \uu2.w_addr_displaying_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4_rep1C_net\,
            ce => 'H',
            sr => \N__15851\
        );

    \uu2.w_addr_displaying_fast_RNILLSO_7_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16458\,
            in1 => \N__14222\,
            in2 => \N__16417\,
            in3 => \N__14790\,
            lcout => \uu2.Z_decfrac106_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_5_rep1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__16463\,
            in1 => \N__13925\,
            in2 => \_gnd_net_\,
            in3 => \N__16055\,
            lcout => \uu2.w_addr_displaying_5_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4_rep1C_net\,
            ce => 'H',
            sr => \N__15851\
        );

    \uu2.w_addr_displaying_fast_7_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100100000"
        )
    port map (
            in0 => \N__16053\,
            in1 => \N__14011\,
            in2 => \N__13929\,
            in3 => \N__14223\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4_rep1C_net\,
            ce => 'H',
            sr => \N__15851\
        );

    \uu2.w_addr_displaying_4_rep1_RNI65VM_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__14820\,
            in1 => \N__15441\,
            in2 => \N__13857\,
            in3 => \N__14890\,
            lcout => \uu2.un1_w_addr_displaying_35_0\,
            ltout => \uu2.un1_w_addr_displaying_35_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIPHFA2_4_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__14461\,
            in1 => \N__13779\,
            in2 => \N__13683\,
            in3 => \N__13679\,
            lcout => \uu2.N_813_0\,
            ltout => \uu2.N_813_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_58_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__16595\,
            in1 => \N__14415\,
            in2 => \N__13668\,
            in3 => \N__14369\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep1_RNIAVDB_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__14891\,
            in1 => \N__14821\,
            in2 => \_gnd_net_\,
            in3 => \N__15442\,
            lcout => \uu2.un1_segment3_m4_s_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec0.segmentUQ_3_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010111101"
        )
    port map (
            in0 => \N__14749\,
            in1 => \N__17239\,
            in2 => \N__14679\,
            in3 => \N__15725\,
            lcout => OPEN,
            ltout => \L3_segment1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIQD7R4_5_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__14580\,
            in1 => \N__14572\,
            in2 => \N__14514\,
            in3 => \N__14503\,
            lcout => \uu2.w_addr_displaying_fast_RNIQD7R4Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIL396_8_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14221\,
            in2 => \N__15240\,
            in3 => \_gnd_net_\,
            lcout => \uu2.N_315_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_59_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111110000"
        )
    port map (
            in0 => \N__14416\,
            in1 => \N__16596\,
            in2 => \N__14384\,
            in3 => \N__14346\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_rep1_RNIUV0B3_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__16252\,
            in1 => \N__14286\,
            in2 => \N__14331\,
            in3 => \N__16491\,
            lcout => \uu2.segment2_m_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_rep1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__14287\,
            in1 => \_gnd_net_\,
            in2 => \N__16095\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displaying_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0_rep1C_net\,
            ce => 'H',
            sr => \N__15856\
        );

    \uu2.w_addr_displaying_4_rep2_RNI4S6J_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__15420\,
            in1 => \N__14284\,
            in2 => \_gnd_net_\,
            in3 => \N__15526\,
            lcout => \uu2.w_addr_displaying_4_rep2_RNI4S6JZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIEDBM_7_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010000000000"
        )
    port map (
            in0 => \N__14285\,
            in1 => \N__15421\,
            in2 => \N__15545\,
            in3 => \N__14233\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_fast_RNIEDBMZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNITRMC1_8_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__15235\,
            in1 => \N__15570\,
            in2 => \N__15564\,
            in3 => \_gnd_net_\,
            lcout => \uu2.un1_segment4_sn_N_38_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep2_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101001101010"
        )
    port map (
            in0 => \N__15530\,
            in1 => \N__15307\,
            in2 => \N__16096\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displaying_4_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0_rep1C_net\,
            ce => 'H',
            sr => \N__15856\
        );

    \uu2.w_addr_displaying_3_rep1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15491\,
            in2 => \N__15449\,
            in3 => \N__16065\,
            lcout => \uu2.w_addr_displaying_3_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0_rep1C_net\,
            ce => 'H',
            sr => \N__15856\
        );

    \uu2.w_addr_displaying_fast_8_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__16066\,
            in1 => \N__15236\,
            in2 => \N__15368\,
            in3 => \N__15308\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0_rep1C_net\,
            ce => 'H',
            sr => \N__15856\
        );

    \Lab_UT.dec3.segmentUQ_2_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__15182\,
            in1 => \N__17050\,
            in2 => \N__15100\,
            in3 => \N__17443\,
            lcout => OPEN,
            ltout => \L3_segment4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_rep1_RNIABAE_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16344\,
            in1 => \_gnd_net_\,
            in2 => \N__15198\,
            in3 => \N__15009\,
            lcout => \uu2.N_280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dec3.segmentUQ_4_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011111101"
        )
    port map (
            in0 => \N__15183\,
            in1 => \N__17049\,
            in2 => \N__15101\,
            in3 => \N__17442\,
            lcout => \L3_segment4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_rep1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__16345\,
            in1 => \N__16136\,
            in2 => \N__16097\,
            in3 => \N__15003\,
            lcout => \uu2.w_addr_displaying_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__15858\
        );

    \uu2.w_addr_displaying_5_rep1_RNI9Q311_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__16465\,
            in1 => \N__16416\,
            in2 => \_gnd_net_\,
            in3 => \N__16342\,
            lcout => \uu2.un1_w_addr_displaying_46_1\,
            ltout => \uu2.un1_w_addr_displaying_46_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI8U3D2_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16135\,
            in2 => \N__16485\,
            in3 => \N__16311\,
            lcout => \uu2.w_addr_displaying_RNI8U3D2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_5_rep1_RNI9Q311_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__16464\,
            in1 => \N__16415\,
            in2 => \_gnd_net_\,
            in3 => \N__16343\,
            lcout => \uu2.un1_w_addr_displaying_38_1\,
            ltout => \uu2.un1_w_addr_displaying_38_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIBSR63_7_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__16305\,
            in1 => \N__16134\,
            in2 => \N__16293\,
            in3 => \N__16253\,
            lcout => \uu2.segment3_m_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16094\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16152\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0C_net\,
            ce => 'H',
            sr => \N__15859\
        );

    \uu2.w_addr_displaying_fast_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16093\,
            in2 => \_gnd_net_\,
            in3 => \N__15943\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0C_net\,
            ce => 'H',
            sr => \N__15859\
        );

    \uu2.mem0.ram512X8_inst_RNO_60_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111111101101"
        )
    port map (
            in0 => \N__16938\,
            in1 => \N__16855\,
            in2 => \N__16681\,
            in3 => \N__16780\,
            lcout => \uu2.mem0.N_2160_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15735\,
            in1 => \N__17112\,
            in2 => \_gnd_net_\,
            in3 => \N__15654\,
            lcout => OPEN,
            ltout => \Lab_UT.didpuu0.ledDisp00.selLed_RNI3BF11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNITQOS1_1_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__17166\,
            in1 => \_gnd_net_\,
            in2 => \N__17466\,
            in3 => \N__17349\,
            lcout => led_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNINURJ_0_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17451\,
            in1 => \N__16669\,
            in2 => \_gnd_net_\,
            in3 => \N__17114\,
            lcout => \Lab_UT.didpuu0.ledDisp00.selLed_RNINURJZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11_0_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17113\,
            in1 => \N__17343\,
            in2 => \_gnd_net_\,
            in3 => \N__17254\,
            lcout => OPEN,
            ltout => \Lab_UT.didpuu0.ledDisp00.selLed_RNI5DF11Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNI1VOS1_1_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__16977\,
            in1 => \_gnd_net_\,
            in2 => \N__17169\,
            in3 => \N__17165\,
            lcout => led_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJ_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__17115\,
            in1 => \_gnd_net_\,
            in2 => \N__16873\,
            in3 => \N__17062\,
            lcout => \Lab_UT.didpuu0.ledDisp00.selLed_RNIP0SJZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.g0_i_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__16932\,
            in1 => \N__16848\,
            in2 => \N__16783\,
            in3 => \N__16661\,
            lcout => \uu2.N_2160_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didpuu0.o_oneSecPluse_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16581\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16548\,
            lcout => led_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

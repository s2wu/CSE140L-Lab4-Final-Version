// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Feb 25 2020 07:08:25

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__13611;
    wire N__13610;
    wire N__13609;
    wire N__13602;
    wire N__13601;
    wire N__13600;
    wire N__13593;
    wire N__13592;
    wire N__13591;
    wire N__13584;
    wire N__13583;
    wire N__13582;
    wire N__13575;
    wire N__13574;
    wire N__13573;
    wire N__13566;
    wire N__13565;
    wire N__13564;
    wire N__13557;
    wire N__13556;
    wire N__13555;
    wire N__13548;
    wire N__13547;
    wire N__13546;
    wire N__13539;
    wire N__13538;
    wire N__13537;
    wire N__13530;
    wire N__13529;
    wire N__13528;
    wire N__13511;
    wire N__13510;
    wire N__13507;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13492;
    wire N__13487;
    wire N__13486;
    wire N__13483;
    wire N__13480;
    wire N__13479;
    wire N__13474;
    wire N__13471;
    wire N__13468;
    wire N__13463;
    wire N__13462;
    wire N__13459;
    wire N__13456;
    wire N__13453;
    wire N__13452;
    wire N__13449;
    wire N__13446;
    wire N__13443;
    wire N__13438;
    wire N__13433;
    wire N__13432;
    wire N__13431;
    wire N__13430;
    wire N__13429;
    wire N__13428;
    wire N__13427;
    wire N__13426;
    wire N__13425;
    wire N__13424;
    wire N__13423;
    wire N__13422;
    wire N__13421;
    wire N__13420;
    wire N__13419;
    wire N__13418;
    wire N__13417;
    wire N__13416;
    wire N__13415;
    wire N__13414;
    wire N__13413;
    wire N__13412;
    wire N__13411;
    wire N__13410;
    wire N__13409;
    wire N__13408;
    wire N__13407;
    wire N__13406;
    wire N__13405;
    wire N__13404;
    wire N__13403;
    wire N__13402;
    wire N__13401;
    wire N__13400;
    wire N__13399;
    wire N__13398;
    wire N__13397;
    wire N__13396;
    wire N__13395;
    wire N__13394;
    wire N__13393;
    wire N__13392;
    wire N__13391;
    wire N__13390;
    wire N__13389;
    wire N__13388;
    wire N__13387;
    wire N__13386;
    wire N__13385;
    wire N__13384;
    wire N__13383;
    wire N__13382;
    wire N__13381;
    wire N__13380;
    wire N__13379;
    wire N__13378;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13255;
    wire N__13252;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13232;
    wire N__13229;
    wire N__13228;
    wire N__13227;
    wire N__13226;
    wire N__13225;
    wire N__13224;
    wire N__13223;
    wire N__13220;
    wire N__13211;
    wire N__13210;
    wire N__13209;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13189;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13161;
    wire N__13160;
    wire N__13155;
    wire N__13150;
    wire N__13145;
    wire N__13144;
    wire N__13141;
    wire N__13140;
    wire N__13137;
    wire N__13136;
    wire N__13131;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13121;
    wire N__13118;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13108;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13094;
    wire N__13091;
    wire N__13086;
    wire N__13083;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13067;
    wire N__13066;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13055;
    wire N__13054;
    wire N__13051;
    wire N__13044;
    wire N__13041;
    wire N__13040;
    wire N__13033;
    wire N__13032;
    wire N__13031;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13017;
    wire N__13010;
    wire N__13007;
    wire N__13004;
    wire N__13001;
    wire N__13000;
    wire N__12999;
    wire N__12998;
    wire N__12995;
    wire N__12992;
    wire N__12991;
    wire N__12988;
    wire N__12985;
    wire N__12984;
    wire N__12983;
    wire N__12980;
    wire N__12979;
    wire N__12976;
    wire N__12967;
    wire N__12966;
    wire N__12963;
    wire N__12962;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12943;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12919;
    wire N__12916;
    wire N__12915;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12903;
    wire N__12900;
    wire N__12895;
    wire N__12892;
    wire N__12889;
    wire N__12886;
    wire N__12881;
    wire N__12880;
    wire N__12877;
    wire N__12876;
    wire N__12875;
    wire N__12874;
    wire N__12873;
    wire N__12872;
    wire N__12871;
    wire N__12868;
    wire N__12867;
    wire N__12864;
    wire N__12861;
    wire N__12860;
    wire N__12857;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12832;
    wire N__12829;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12808;
    wire N__12805;
    wire N__12804;
    wire N__12803;
    wire N__12802;
    wire N__12799;
    wire N__12798;
    wire N__12797;
    wire N__12796;
    wire N__12793;
    wire N__12792;
    wire N__12791;
    wire N__12788;
    wire N__12787;
    wire N__12784;
    wire N__12777;
    wire N__12774;
    wire N__12773;
    wire N__12770;
    wire N__12769;
    wire N__12766;
    wire N__12763;
    wire N__12760;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12748;
    wire N__12739;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12719;
    wire N__12710;
    wire N__12707;
    wire N__12706;
    wire N__12705;
    wire N__12702;
    wire N__12699;
    wire N__12698;
    wire N__12695;
    wire N__12694;
    wire N__12693;
    wire N__12692;
    wire N__12687;
    wire N__12686;
    wire N__12685;
    wire N__12684;
    wire N__12683;
    wire N__12682;
    wire N__12681;
    wire N__12678;
    wire N__12677;
    wire N__12676;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12651;
    wire N__12644;
    wire N__12637;
    wire N__12634;
    wire N__12629;
    wire N__12614;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12602;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12598;
    wire N__12595;
    wire N__12592;
    wire N__12591;
    wire N__12590;
    wire N__12587;
    wire N__12586;
    wire N__12585;
    wire N__12584;
    wire N__12581;
    wire N__12576;
    wire N__12567;
    wire N__12564;
    wire N__12563;
    wire N__12562;
    wire N__12561;
    wire N__12558;
    wire N__12555;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12541;
    wire N__12538;
    wire N__12533;
    wire N__12530;
    wire N__12525;
    wire N__12522;
    wire N__12509;
    wire N__12508;
    wire N__12505;
    wire N__12504;
    wire N__12503;
    wire N__12502;
    wire N__12501;
    wire N__12500;
    wire N__12499;
    wire N__12498;
    wire N__12497;
    wire N__12496;
    wire N__12495;
    wire N__12494;
    wire N__12493;
    wire N__12490;
    wire N__12489;
    wire N__12488;
    wire N__12487;
    wire N__12486;
    wire N__12485;
    wire N__12476;
    wire N__12469;
    wire N__12468;
    wire N__12467;
    wire N__12466;
    wire N__12465;
    wire N__12464;
    wire N__12463;
    wire N__12462;
    wire N__12457;
    wire N__12450;
    wire N__12447;
    wire N__12442;
    wire N__12433;
    wire N__12428;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12394;
    wire N__12377;
    wire N__12374;
    wire N__12371;
    wire N__12370;
    wire N__12367;
    wire N__12362;
    wire N__12359;
    wire N__12358;
    wire N__12357;
    wire N__12356;
    wire N__12355;
    wire N__12352;
    wire N__12349;
    wire N__12346;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12332;
    wire N__12323;
    wire N__12322;
    wire N__12321;
    wire N__12318;
    wire N__12313;
    wire N__12312;
    wire N__12311;
    wire N__12310;
    wire N__12309;
    wire N__12308;
    wire N__12307;
    wire N__12306;
    wire N__12305;
    wire N__12304;
    wire N__12303;
    wire N__12302;
    wire N__12301;
    wire N__12300;
    wire N__12299;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12291;
    wire N__12290;
    wire N__12289;
    wire N__12288;
    wire N__12287;
    wire N__12286;
    wire N__12285;
    wire N__12284;
    wire N__12283;
    wire N__12282;
    wire N__12281;
    wire N__12224;
    wire N__12221;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12202;
    wire N__12199;
    wire N__12196;
    wire N__12191;
    wire N__12188;
    wire N__12187;
    wire N__12186;
    wire N__12183;
    wire N__12178;
    wire N__12173;
    wire N__12172;
    wire N__12169;
    wire N__12168;
    wire N__12165;
    wire N__12162;
    wire N__12159;
    wire N__12156;
    wire N__12151;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12137;
    wire N__12136;
    wire N__12133;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12121;
    wire N__12116;
    wire N__12113;
    wire N__12112;
    wire N__12111;
    wire N__12108;
    wire N__12103;
    wire N__12098;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12079;
    wire N__12078;
    wire N__12077;
    wire N__12074;
    wire N__12073;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12065;
    wire N__12064;
    wire N__12063;
    wire N__12060;
    wire N__12059;
    wire N__12056;
    wire N__12051;
    wire N__12050;
    wire N__12049;
    wire N__12046;
    wire N__12043;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12029;
    wire N__12024;
    wire N__12019;
    wire N__12012;
    wire N__11999;
    wire N__11996;
    wire N__11993;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11983;
    wire N__11982;
    wire N__11979;
    wire N__11974;
    wire N__11971;
    wire N__11968;
    wire N__11967;
    wire N__11966;
    wire N__11963;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11945;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11935;
    wire N__11934;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11924;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11906;
    wire N__11905;
    wire N__11900;
    wire N__11899;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11872;
    wire N__11869;
    wire N__11866;
    wire N__11865;
    wire N__11864;
    wire N__11863;
    wire N__11860;
    wire N__11857;
    wire N__11852;
    wire N__11849;
    wire N__11848;
    wire N__11847;
    wire N__11840;
    wire N__11835;
    wire N__11832;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11818;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11803;
    wire N__11800;
    wire N__11795;
    wire N__11794;
    wire N__11791;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11735;
    wire N__11732;
    wire N__11731;
    wire N__11730;
    wire N__11729;
    wire N__11726;
    wire N__11721;
    wire N__11720;
    wire N__11719;
    wire N__11716;
    wire N__11711;
    wire N__11704;
    wire N__11699;
    wire N__11696;
    wire N__11695;
    wire N__11694;
    wire N__11693;
    wire N__11692;
    wire N__11687;
    wire N__11684;
    wire N__11683;
    wire N__11678;
    wire N__11677;
    wire N__11676;
    wire N__11675;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11653;
    wire N__11646;
    wire N__11639;
    wire N__11638;
    wire N__11637;
    wire N__11634;
    wire N__11633;
    wire N__11630;
    wire N__11629;
    wire N__11628;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11609;
    wire N__11606;
    wire N__11597;
    wire N__11596;
    wire N__11593;
    wire N__11592;
    wire N__11591;
    wire N__11590;
    wire N__11587;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11575;
    wire N__11572;
    wire N__11571;
    wire N__11568;
    wire N__11565;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11547;
    wire N__11544;
    wire N__11531;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11502;
    wire N__11497;
    wire N__11494;
    wire N__11489;
    wire N__11488;
    wire N__11487;
    wire N__11484;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11476;
    wire N__11465;
    wire N__11462;
    wire N__11459;
    wire N__11458;
    wire N__11457;
    wire N__11456;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11448;
    wire N__11445;
    wire N__11440;
    wire N__11437;
    wire N__11432;
    wire N__11427;
    wire N__11420;
    wire N__11417;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11409;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11387;
    wire N__11386;
    wire N__11383;
    wire N__11382;
    wire N__11379;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11357;
    wire N__11356;
    wire N__11355;
    wire N__11354;
    wire N__11351;
    wire N__11344;
    wire N__11343;
    wire N__11338;
    wire N__11335;
    wire N__11330;
    wire N__11329;
    wire N__11324;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11299;
    wire N__11298;
    wire N__11295;
    wire N__11290;
    wire N__11285;
    wire N__11284;
    wire N__11281;
    wire N__11280;
    wire N__11279;
    wire N__11278;
    wire N__11277;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11259;
    wire N__11252;
    wire N__11251;
    wire N__11250;
    wire N__11249;
    wire N__11248;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11244;
    wire N__11243;
    wire N__11242;
    wire N__11237;
    wire N__11224;
    wire N__11221;
    wire N__11220;
    wire N__11219;
    wire N__11218;
    wire N__11217;
    wire N__11214;
    wire N__11213;
    wire N__11210;
    wire N__11205;
    wire N__11202;
    wire N__11201;
    wire N__11198;
    wire N__11193;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11183;
    wire N__11180;
    wire N__11175;
    wire N__11172;
    wire N__11169;
    wire N__11166;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11150;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11113;
    wire N__11110;
    wire N__11107;
    wire N__11102;
    wire N__11101;
    wire N__11096;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11088;
    wire N__11087;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11073;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11046;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11023;
    wire N__11020;
    wire N__11017;
    wire N__11012;
    wire N__11009;
    wire N__11008;
    wire N__11007;
    wire N__11006;
    wire N__11005;
    wire N__11002;
    wire N__10993;
    wire N__10988;
    wire N__10987;
    wire N__10986;
    wire N__10985;
    wire N__10984;
    wire N__10981;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10942;
    wire N__10937;
    wire N__10936;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10925;
    wire N__10924;
    wire N__10921;
    wire N__10920;
    wire N__10919;
    wire N__10918;
    wire N__10917;
    wire N__10916;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10902;
    wire N__10895;
    wire N__10890;
    wire N__10885;
    wire N__10874;
    wire N__10873;
    wire N__10872;
    wire N__10869;
    wire N__10868;
    wire N__10867;
    wire N__10864;
    wire N__10863;
    wire N__10860;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10840;
    wire N__10829;
    wire N__10826;
    wire N__10825;
    wire N__10822;
    wire N__10821;
    wire N__10820;
    wire N__10819;
    wire N__10818;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10799;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10783;
    wire N__10782;
    wire N__10779;
    wire N__10774;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10762;
    wire N__10761;
    wire N__10760;
    wire N__10755;
    wire N__10754;
    wire N__10753;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10735;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10696;
    wire N__10695;
    wire N__10692;
    wire N__10691;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10679;
    wire N__10676;
    wire N__10675;
    wire N__10674;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10666;
    wire N__10665;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10650;
    wire N__10645;
    wire N__10638;
    wire N__10625;
    wire N__10624;
    wire N__10621;
    wire N__10620;
    wire N__10619;
    wire N__10618;
    wire N__10617;
    wire N__10614;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10596;
    wire N__10595;
    wire N__10592;
    wire N__10591;
    wire N__10588;
    wire N__10583;
    wire N__10580;
    wire N__10579;
    wire N__10578;
    wire N__10575;
    wire N__10568;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10519;
    wire N__10518;
    wire N__10517;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10509;
    wire N__10508;
    wire N__10507;
    wire N__10506;
    wire N__10505;
    wire N__10500;
    wire N__10497;
    wire N__10494;
    wire N__10489;
    wire N__10488;
    wire N__10487;
    wire N__10486;
    wire N__10485;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10477;
    wire N__10476;
    wire N__10473;
    wire N__10472;
    wire N__10471;
    wire N__10470;
    wire N__10469;
    wire N__10466;
    wire N__10457;
    wire N__10450;
    wire N__10445;
    wire N__10438;
    wire N__10431;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10393;
    wire N__10390;
    wire N__10389;
    wire N__10384;
    wire N__10381;
    wire N__10376;
    wire N__10373;
    wire N__10372;
    wire N__10371;
    wire N__10368;
    wire N__10367;
    wire N__10362;
    wire N__10357;
    wire N__10352;
    wire N__10349;
    wire N__10348;
    wire N__10347;
    wire N__10344;
    wire N__10339;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10324;
    wire N__10323;
    wire N__10322;
    wire N__10321;
    wire N__10320;
    wire N__10319;
    wire N__10318;
    wire N__10317;
    wire N__10310;
    wire N__10303;
    wire N__10296;
    wire N__10289;
    wire N__10288;
    wire N__10287;
    wire N__10286;
    wire N__10285;
    wire N__10284;
    wire N__10281;
    wire N__10280;
    wire N__10279;
    wire N__10278;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10274;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10254;
    wire N__10245;
    wire N__10244;
    wire N__10241;
    wire N__10240;
    wire N__10239;
    wire N__10238;
    wire N__10237;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10223;
    wire N__10216;
    wire N__10207;
    wire N__10204;
    wire N__10193;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10159;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10144;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10096;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10082;
    wire N__10079;
    wire N__10078;
    wire N__10077;
    wire N__10076;
    wire N__10069;
    wire N__10066;
    wire N__10065;
    wire N__10060;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10050;
    wire N__10047;
    wire N__10044;
    wire N__10039;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10018;
    wire N__10015;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__10007;
    wire N__10006;
    wire N__10005;
    wire N__10002;
    wire N__9999;
    wire N__9996;
    wire N__9989;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9967;
    wire N__9966;
    wire N__9965;
    wire N__9964;
    wire N__9961;
    wire N__9958;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9946;
    wire N__9945;
    wire N__9944;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9929;
    wire N__9922;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9902;
    wire N__9901;
    wire N__9900;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9888;
    wire N__9885;
    wire N__9880;
    wire N__9875;
    wire N__9872;
    wire N__9871;
    wire N__9870;
    wire N__9869;
    wire N__9866;
    wire N__9865;
    wire N__9862;
    wire N__9861;
    wire N__9858;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9844;
    wire N__9843;
    wire N__9842;
    wire N__9839;
    wire N__9834;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9800;
    wire N__9797;
    wire N__9796;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9788;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9773;
    wire N__9764;
    wire N__9763;
    wire N__9762;
    wire N__9761;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9750;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9738;
    wire N__9731;
    wire N__9726;
    wire N__9723;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9707;
    wire N__9706;
    wire N__9705;
    wire N__9704;
    wire N__9703;
    wire N__9700;
    wire N__9699;
    wire N__9696;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9672;
    wire N__9671;
    wire N__9670;
    wire N__9669;
    wire N__9664;
    wire N__9659;
    wire N__9654;
    wire N__9649;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9617;
    wire N__9616;
    wire N__9615;
    wire N__9608;
    wire N__9605;
    wire N__9604;
    wire N__9603;
    wire N__9602;
    wire N__9599;
    wire N__9598;
    wire N__9597;
    wire N__9590;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9582;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9556;
    wire N__9545;
    wire N__9544;
    wire N__9541;
    wire N__9540;
    wire N__9539;
    wire N__9538;
    wire N__9535;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9527;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9513;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9497;
    wire N__9494;
    wire N__9489;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9463;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9448;
    wire N__9445;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9421;
    wire N__9420;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9412;
    wire N__9411;
    wire N__9410;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9371;
    wire N__9370;
    wire N__9369;
    wire N__9362;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9344;
    wire N__9343;
    wire N__9342;
    wire N__9339;
    wire N__9338;
    wire N__9331;
    wire N__9328;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9313;
    wire N__9312;
    wire N__9311;
    wire N__9308;
    wire N__9301;
    wire N__9296;
    wire N__9293;
    wire N__9292;
    wire N__9291;
    wire N__9290;
    wire N__9281;
    wire N__9280;
    wire N__9279;
    wire N__9276;
    wire N__9273;
    wire N__9270;
    wire N__9267;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9238;
    wire N__9237;
    wire N__9236;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9228;
    wire N__9225;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9210;
    wire N__9209;
    wire N__9206;
    wire N__9205;
    wire N__9204;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9188;
    wire N__9185;
    wire N__9180;
    wire N__9167;
    wire N__9164;
    wire N__9163;
    wire N__9162;
    wire N__9157;
    wire N__9156;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9138;
    wire N__9137;
    wire N__9136;
    wire N__9135;
    wire N__9134;
    wire N__9133;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9110;
    wire N__9103;
    wire N__9100;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9052;
    wire N__9051;
    wire N__9050;
    wire N__9047;
    wire N__9040;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9007;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8999;
    wire N__8996;
    wire N__8989;
    wire N__8984;
    wire N__8983;
    wire N__8982;
    wire N__8981;
    wire N__8980;
    wire N__8975;
    wire N__8968;
    wire N__8963;
    wire N__8960;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8893;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8866;
    wire N__8863;
    wire N__8858;
    wire N__8855;
    wire N__8854;
    wire N__8853;
    wire N__8848;
    wire N__8847;
    wire N__8846;
    wire N__8845;
    wire N__8844;
    wire N__8843;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8829;
    wire N__8822;
    wire N__8819;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8785;
    wire N__8782;
    wire N__8781;
    wire N__8778;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8755;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8704;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8692;
    wire N__8687;
    wire N__8684;
    wire N__8683;
    wire N__8680;
    wire N__8677;
    wire N__8674;
    wire N__8669;
    wire N__8668;
    wire N__8663;
    wire N__8660;
    wire N__8659;
    wire N__8656;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8639;
    wire N__8638;
    wire N__8637;
    wire N__8636;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8618;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8584;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8549;
    wire N__8548;
    wire N__8547;
    wire N__8546;
    wire N__8543;
    wire N__8538;
    wire N__8535;
    wire N__8534;
    wire N__8529;
    wire N__8526;
    wire N__8525;
    wire N__8522;
    wire N__8521;
    wire N__8520;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8506;
    wire N__8503;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8473;
    wire N__8468;
    wire N__8467;
    wire N__8466;
    wire N__8463;
    wire N__8462;
    wire N__8461;
    wire N__8456;
    wire N__8453;
    wire N__8448;
    wire N__8441;
    wire N__8438;
    wire N__8437;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8409;
    wire N__8408;
    wire N__8407;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8399;
    wire N__8398;
    wire N__8397;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8366;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8332;
    wire N__8329;
    wire N__8328;
    wire N__8325;
    wire N__8324;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8314;
    wire N__8313;
    wire N__8312;
    wire N__8311;
    wire N__8310;
    wire N__8309;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8297;
    wire N__8292;
    wire N__8287;
    wire N__8280;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8251;
    wire N__8250;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8230;
    wire N__8229;
    wire N__8224;
    wire N__8221;
    wire N__8216;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8206;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8179;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8167;
    wire N__8166;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8141;
    wire N__8140;
    wire N__8139;
    wire N__8138;
    wire N__8137;
    wire N__8128;
    wire N__8125;
    wire N__8120;
    wire N__8119;
    wire N__8116;
    wire N__8115;
    wire N__8112;
    wire N__8111;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8097;
    wire N__8092;
    wire N__8087;
    wire N__8086;
    wire N__8085;
    wire N__8082;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8061;
    wire N__8058;
    wire N__8055;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8032;
    wire N__8031;
    wire N__8028;
    wire N__8025;
    wire N__8022;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__7997;
    wire N__7996;
    wire N__7991;
    wire N__7988;
    wire N__7987;
    wire N__7986;
    wire N__7985;
    wire N__7982;
    wire N__7975;
    wire N__7970;
    wire N__7969;
    wire N__7968;
    wire N__7967;
    wire N__7966;
    wire N__7963;
    wire N__7954;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7930;
    wire N__7929;
    wire N__7928;
    wire N__7927;
    wire N__7924;
    wire N__7923;
    wire N__7914;
    wire N__7911;
    wire N__7908;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7876;
    wire N__7875;
    wire N__7870;
    wire N__7867;
    wire N__7864;
    wire N__7859;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7804;
    wire N__7803;
    wire N__7800;
    wire N__7799;
    wire N__7796;
    wire N__7793;
    wire N__7792;
    wire N__7789;
    wire N__7780;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7741;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7657;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7558;
    wire N__7557;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7541;
    wire N__7538;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7514;
    wire N__7513;
    wire N__7512;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7500;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7474;
    wire N__7471;
    wire N__7470;
    wire N__7469;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7455;
    wire N__7454;
    wire N__7453;
    wire N__7446;
    wire N__7445;
    wire N__7444;
    wire N__7443;
    wire N__7442;
    wire N__7437;
    wire N__7434;
    wire N__7425;
    wire N__7418;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7410;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7398;
    wire N__7391;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7300;
    wire N__7297;
    wire N__7296;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7282;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7268;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7250;
    wire N__7247;
    wire N__7246;
    wire N__7243;
    wire N__7240;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7190;
    wire N__7187;
    wire N__7184;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7156;
    wire N__7155;
    wire N__7152;
    wire N__7147;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7003;
    wire N__6998;
    wire N__6995;
    wire N__6992;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6980;
    wire N__6977;
    wire N__6976;
    wire N__6975;
    wire N__6970;
    wire N__6967;
    wire N__6962;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6952;
    wire N__6949;
    wire N__6944;
    wire N__6943;
    wire N__6942;
    wire N__6939;
    wire N__6934;
    wire N__6929;
    wire N__6926;
    wire N__6925;
    wire N__6924;
    wire N__6923;
    wire N__6920;
    wire N__6913;
    wire N__6910;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6802;
    wire N__6801;
    wire N__6800;
    wire N__6791;
    wire N__6788;
    wire N__6787;
    wire N__6786;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6772;
    wire N__6769;
    wire N__6766;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6754;
    wire N__6753;
    wire N__6752;
    wire N__6743;
    wire N__6740;
    wire N__6739;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6727;
    wire N__6724;
    wire N__6723;
    wire N__6720;
    wire N__6719;
    wire N__6718;
    wire N__6717;
    wire N__6714;
    wire N__6713;
    wire N__6710;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6667;
    wire N__6666;
    wire N__6661;
    wire N__6658;
    wire N__6653;
    wire N__6652;
    wire N__6651;
    wire N__6650;
    wire N__6643;
    wire N__6640;
    wire N__6635;
    wire N__6634;
    wire N__6633;
    wire N__6632;
    wire N__6629;
    wire N__6628;
    wire N__6625;
    wire N__6618;
    wire N__6615;
    wire N__6608;
    wire N__6607;
    wire N__6606;
    wire N__6605;
    wire N__6602;
    wire N__6595;
    wire N__6592;
    wire N__6587;
    wire N__6584;
    wire N__6583;
    wire N__6582;
    wire N__6581;
    wire N__6578;
    wire N__6577;
    wire N__6576;
    wire N__6575;
    wire N__6574;
    wire N__6573;
    wire N__6572;
    wire N__6569;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6557;
    wire N__6546;
    wire N__6541;
    wire N__6530;
    wire N__6529;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6517;
    wire N__6514;
    wire N__6513;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6501;
    wire N__6498;
    wire N__6491;
    wire N__6488;
    wire N__6487;
    wire N__6486;
    wire N__6485;
    wire N__6484;
    wire N__6483;
    wire N__6482;
    wire N__6477;
    wire N__6472;
    wire N__6465;
    wire N__6464;
    wire N__6463;
    wire N__6462;
    wire N__6461;
    wire N__6460;
    wire N__6453;
    wire N__6450;
    wire N__6441;
    wire N__6434;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6421;
    wire N__6418;
    wire N__6417;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6402;
    wire N__6395;
    wire N__6392;
    wire N__6391;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6374;
    wire N__6373;
    wire N__6372;
    wire N__6371;
    wire N__6370;
    wire N__6359;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6286;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6269;
    wire N__6268;
    wire N__6267;
    wire N__6264;
    wire N__6257;
    wire N__6254;
    wire N__6253;
    wire N__6252;
    wire N__6251;
    wire N__6248;
    wire N__6241;
    wire N__6238;
    wire N__6233;
    wire N__6230;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6218;
    wire N__6217;
    wire N__6214;
    wire N__6213;
    wire N__6212;
    wire N__6209;
    wire N__6208;
    wire N__6205;
    wire N__6198;
    wire N__6195;
    wire N__6188;
    wire N__6187;
    wire N__6186;
    wire N__6183;
    wire N__6176;
    wire N__6173;
    wire N__6172;
    wire N__6169;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6159;
    wire N__6152;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6140;
    wire N__6137;
    wire N__6136;
    wire N__6135;
    wire N__6134;
    wire N__6131;
    wire N__6124;
    wire N__6121;
    wire N__6116;
    wire N__6113;
    wire N__6112;
    wire N__6111;
    wire N__6106;
    wire N__6103;
    wire N__6098;
    wire N__6097;
    wire N__6094;
    wire N__6093;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6081;
    wire N__6078;
    wire N__6071;
    wire N__6068;
    wire N__6067;
    wire N__6066;
    wire N__6065;
    wire N__6064;
    wire N__6061;
    wire N__6054;
    wire N__6051;
    wire N__6044;
    wire N__6043;
    wire N__6040;
    wire N__6039;
    wire N__6038;
    wire N__6037;
    wire N__6036;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6016;
    wire N__6015;
    wire N__6014;
    wire N__6013;
    wire N__6010;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5988;
    wire N__5983;
    wire N__5978;
    wire N__5977;
    wire N__5976;
    wire N__5975;
    wire N__5972;
    wire N__5965;
    wire N__5962;
    wire N__5957;
    wire N__5956;
    wire N__5955;
    wire N__5954;
    wire N__5953;
    wire N__5944;
    wire N__5941;
    wire N__5936;
    wire N__5935;
    wire N__5932;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5917;
    wire N__5912;
    wire N__5911;
    wire N__5910;
    wire N__5907;
    wire N__5902;
    wire N__5899;
    wire N__5894;
    wire N__5893;
    wire N__5892;
    wire N__5887;
    wire N__5884;
    wire N__5879;
    wire N__5876;
    wire N__5875;
    wire N__5874;
    wire N__5873;
    wire N__5872;
    wire N__5863;
    wire N__5860;
    wire N__5855;
    wire N__5852;
    wire N__5851;
    wire N__5850;
    wire N__5847;
    wire N__5842;
    wire N__5839;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5817;
    wire N__5816;
    wire N__5815;
    wire N__5814;
    wire N__5813;
    wire N__5812;
    wire N__5809;
    wire N__5806;
    wire N__5793;
    wire N__5788;
    wire N__5785;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5773;
    wire N__5772;
    wire N__5769;
    wire N__5768;
    wire N__5761;
    wire N__5758;
    wire N__5753;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5745;
    wire N__5744;
    wire N__5743;
    wire N__5742;
    wire N__5739;
    wire N__5730;
    wire N__5727;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5671;
    wire N__5668;
    wire N__5667;
    wire N__5664;
    wire N__5663;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5651;
    wire N__5648;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5632;
    wire N__5631;
    wire N__5630;
    wire N__5627;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5609;
    wire N__5608;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5595;
    wire N__5592;
    wire N__5589;
    wire N__5586;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5572;
    wire N__5569;
    wire N__5568;
    wire N__5567;
    wire N__5566;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5549;
    wire N__5546;
    wire N__5537;
    wire N__5536;
    wire N__5535;
    wire N__5534;
    wire N__5533;
    wire N__5526;
    wire N__5521;
    wire N__5518;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5495;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5487;
    wire N__5486;
    wire N__5483;
    wire N__5476;
    wire N__5471;
    wire N__5468;
    wire N__5467;
    wire N__5466;
    wire N__5463;
    wire N__5458;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5446;
    wire N__5445;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5423;
    wire N__5420;
    wire N__5419;
    wire N__5416;
    wire N__5415;
    wire N__5412;
    wire N__5411;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5397;
    wire N__5390;
    wire N__5387;
    wire N__5386;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5338;
    wire N__5333;
    wire N__5330;
    wire N__5329;
    wire N__5328;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5306;
    wire N__5305;
    wire N__5304;
    wire N__5303;
    wire N__5302;
    wire N__5301;
    wire N__5294;
    wire N__5287;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5224;
    wire N__5223;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5215;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5197;
    wire N__5194;
    wire N__5189;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5181;
    wire N__5178;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5156;
    wire N__5153;
    wire N__5152;
    wire N__5151;
    wire N__5146;
    wire N__5143;
    wire N__5138;
    wire N__5135;
    wire N__5134;
    wire N__5133;
    wire N__5132;
    wire N__5129;
    wire N__5124;
    wire N__5119;
    wire N__5114;
    wire N__5113;
    wire N__5112;
    wire N__5111;
    wire N__5106;
    wire N__5101;
    wire N__5096;
    wire N__5093;
    wire N__5092;
    wire N__5091;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire clk_in_c;
    wire GNDG0;
    wire VCCG0;
    wire \resetGen.rst_isoZ0 ;
    wire \Lab_UT.secuu0.un131_ci_3_cascade_ ;
    wire uart_RXD;
    wire \Lab_UT.secuu0.un197_ci_9_cascade_ ;
    wire \Lab_UT.secuu0.un230_ci_1_cascade_ ;
    wire \Lab_UT.secuu0.l_precountZ0Z_0 ;
    wire \Lab_UT.secuu0.l_countZ0Z_4 ;
    wire \Lab_UT.secuu0.un4_l_count_14_cascade_ ;
    wire \Lab_UT.secuu0.un4_l_count_0_8 ;
    wire \Lab_UT.secuu0.un4_l_count_0_8_cascade_ ;
    wire \Lab_UT.secuu0.l_countZ0Z_14 ;
    wire \Lab_UT.secuu0.un197_ci_9 ;
    wire \Lab_UT.secuu0.l_countZ0Z_12 ;
    wire \Lab_UT.secuu0.un208_ci_0 ;
    wire \Lab_UT.secuu0.l_countZ0Z_13 ;
    wire \Lab_UT.secuu0.l_countZ0Z_10 ;
    wire \Lab_UT.secuu0.l_countZ0Z_8 ;
    wire \uu2.mem0.w_addr_8 ;
    wire \uu2.mem0.w_addr_1 ;
    wire \uu2.mem0.w_addr_2 ;
    wire \uu2.mem0.w_addr_5 ;
    wire \uu2.mem0.w_data_4 ;
    wire \uu2.mem0.w_addr_3 ;
    wire \uu2.mem0.g0_0_a3_3_cascade_ ;
    wire \uu2.mem0.w_data_1 ;
    wire \uu2.mem0.g1_0_6_cascade_ ;
    wire \uu2.mem0.N_4_i ;
    wire \uu2.mem0.w_addr_6 ;
    wire \uu2.mem0.N_14_0 ;
    wire \uu2.vbuf_raddr.un459_ci_0_cascade_ ;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.r_addrZ0Z_5 ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \uu2.vbuf_raddr.un437_ci_3 ;
    wire \uu2.un306_ci_cascade_ ;
    wire \uu2.un339_ci_0 ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \uu2.r_addrZ0Z_2 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.r_addrZ0Z_0 ;
    wire \uu2.un415_ci_0 ;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu2.un3_r_clk_en_6_cascade_ ;
    wire uu2_un3_r_clk_en_0_cascade_;
    wire \uu2.vbuf_tx_data_rdy ;
    wire \uu2.un3_r_clk_en_0_0 ;
    wire \uu2.l_countZ0Z_2 ;
    wire \uu2.l_countZ0Z_0 ;
    wire \uu2.un3_r_clk_en_7 ;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \uu2.un372_ci_cascade_ ;
    wire \uu2.l_countZ0Z_10 ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.vbuf_count.un372_ci_8_1 ;
    wire \uu2.l_countZ0Z_8 ;
    wire \uu2.vbuf_count.un372_ci_8_1_cascade_ ;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu2.l_countZ0Z_5 ;
    wire \uu2.un306_ci ;
    wire \uu2.l_countZ0Z_4 ;
    wire \Lab_UT.secuu0.l_precountZ0Z_2 ;
    wire \Lab_UT.secuu0.l_precountZ0Z_1 ;
    wire \Lab_UT.secuu0.l_countZ0Z_5 ;
    wire \Lab_UT.secuu0.l_precountZ0Z_3 ;
    wire \Lab_UT.secuu0.l_countZ0Z_15 ;
    wire \Lab_UT.secuu0.un4_l_count_11_cascade_ ;
    wire \Lab_UT.secuu0.un4_l_count_13 ;
    wire \Lab_UT.secuu0.un4_l_count_16_cascade_ ;
    wire \Lab_UT.secuu0.un4_l_count_18 ;
    wire \Lab_UT.secuu0.delay_lineZ0Z_1 ;
    wire \Lab_UT.secuu0.un4_l_count_0_cascade_ ;
    wire \Lab_UT.secuu0.delay_lineZ0Z_0 ;
    wire \Lab_UT.secuu0.un11_l_count_i ;
    wire \Lab_UT.secuu0.un186_ci_0 ;
    wire \Lab_UT.secuu0.l_countZ0Z_11 ;
    wire \Lab_UT.secuu0.un241_ci_2 ;
    wire \Lab_UT.secuu0.l_countZ0Z_16 ;
    wire \Lab_UT.secuu0.un263_ci_cascade_ ;
    wire \Lab_UT.secuu0.l_countZ0Z_18 ;
    wire \Lab_UT.secuu0.l_countZ0Z_9 ;
    wire \Lab_UT.secuu0.l_countZ0Z_17 ;
    wire \Lab_UT.secuu0.un4_l_count_12 ;
    wire \Lab_UT.secuu0.un87_ci ;
    wire \Lab_UT.secuu0.un87_ci_cascade_ ;
    wire \Lab_UT.secuu0.l_countZ0Z_3 ;
    wire \Lab_UT.secuu0.l_countZ0Z_2 ;
    wire \Lab_UT.secuu0.l_countZ0Z_0 ;
    wire \Lab_UT.secuu0.l_countZ0Z_1 ;
    wire \Lab_UT.secuu0.un109_ci_cascade_ ;
    wire \Lab_UT.secuu0.un153_ci ;
    wire \Lab_UT.secuu0.un131_ci_3 ;
    wire \Lab_UT.secuu0.l_countZ0Z_6 ;
    wire \Lab_UT.secuu0.un4_l_count_0 ;
    wire \Lab_UT.secuu0.un142_ci_0 ;
    wire \Lab_UT.secuu0.un109_ci ;
    wire \Lab_UT.secuu0.l_countZ0Z_7 ;
    wire \Lab_UT.secuu0.un11_l_count_i_g ;
    wire \resetGen.N_104_cascade_ ;
    wire \resetGen.N_84 ;
    wire \resetGen.reset_countZ0Z_0 ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire \resetGen.N_86 ;
    wire \resetGen.N_104 ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire \resetGen.N_86_cascade_ ;
    wire \resetGen.reset_countZ0Z_4 ;
    wire \uu2.mem0.g2_1_0_0_cascade_ ;
    wire \uu2.mem0.g0_2_1 ;
    wire \uu2.mem0.g0_i_a2_3_cascade_ ;
    wire \uu2.mem0.w_data_displaying_2_0_0 ;
    wire \uu2.mem0.g1_0_5 ;
    wire \uu2.mem0.N_10_0_0 ;
    wire \uu2.mem0.g1_2 ;
    wire \uu2.mem0.g1_1_sx ;
    wire \uu2.mem0.g1_0 ;
    wire \uu2.mem0.g0_i_5 ;
    wire \uu2.mem0.g0_i_6_1_0 ;
    wire \uu2.mem0.N_19_cascade_ ;
    wire \uu2.mem0.g0_i_6 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_53 ;
    wire bfn_5_10_0_;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \uu2.mem0.g0_0_a3_0 ;
    wire \buart.Z_rx.startbit_cascade_ ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_rx.ser_clk_cascade_ ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \uu2.r_data_wire_0 ;
    wire \uu2.r_data_wire_1 ;
    wire \uu2.r_data_wire_2 ;
    wire \uu2.r_data_wire_3 ;
    wire \uu2.r_data_wire_4 ;
    wire \uu2.r_data_wire_5 ;
    wire vbuf_tx_data_5;
    wire \uu2.r_data_wire_6 ;
    wire vbuf_tx_data_6;
    wire \uu2.r_data_wire_7 ;
    wire vbuf_tx_data_7;
    wire \uu2.vbuf_tx_data_rdy_0 ;
    wire vbuf_tx_data_3;
    wire vbuf_tx_data_4;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire vbuf_tx_data_2;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire bfn_6_5_0_;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \uu2.mem0.w_data_7 ;
    wire \buart.Z_rx.ser_clk ;
    wire \buart.Z_rx.N_103_cascade_ ;
    wire \resetGen.un3_reset_count_i_a3Z0Z_7 ;
    wire \buart.Z_rx.bitcountZ0Z_4 ;
    wire N_87_cascade_;
    wire \buart.Z_rx.N_91 ;
    wire \buart.Z_rx.N_91_cascade_ ;
    wire \buart.Z_rx.N_29_0_i_2 ;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.N_29_0_i_2_cascade_ ;
    wire \buart.Z_rx.startbit ;
    wire \buart.Z_rx.bitcountZ0Z_1 ;
    wire \buart.Z_rx.bitcounte_0_i_2 ;
    wire \uu2.Z_decfrac105_7_3_cascade_ ;
    wire \uu2.mem0.w_data_6 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_17_cascade_ ;
    wire \uu2.mem0.w_data_5 ;
    wire \uu2.Z_decfrac105_7_3 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_ ;
    wire \uu2.mem0.w_data_0 ;
    wire \INVuu2.w_addr_displaying_5C_net ;
    wire \uu2.mem0.w_data_2 ;
    wire \uu2.un1_w_user_cr_0_0 ;
    wire latticehx1k_pll_inst_PLLOUTCORE_i;
    wire \uu2.un1_w_user_cr_0_0_cascade_ ;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_34_cascade_ ;
    wire \uu2.mem0.un1_segment3_m6_0_0_0_0_cascade_ ;
    wire \uu2.mem0.w_data_3 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_35 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_21 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_22 ;
    wire \uu2.mem0.g0_i_a2_4 ;
    wire \uu2.mem0.N_8_tz_0_0_1 ;
    wire led_c_0_4_cascade_;
    wire \uu2.mem0.g1_0_0_0 ;
    wire \uu2.mem0.g0_i_5_1_0 ;
    wire \uu2.mem0.g2_0 ;
    wire \uu2.w_addr_displaying_4_rep1_8_cascade_ ;
    wire \uu2.N_42_0_0_cascade_ ;
    wire \uu2.N_1482_0_0 ;
    wire \INVuu2.w_addr_displaying_8_rep1C_net ;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire vbuf_tx_data_0;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire vbuf_tx_data_1;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire \uu2.o_adder_vbuf_w_addr_user_3_cascade_ ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.w_addr_userZ1Z_1 ;
    wire \INVuu2.w_addr_user_2C_net ;
    wire \uu2.o_adder_vbuf_w_addr_user_7_cascade_ ;
    wire \uu2.mem0.w_addr_7 ;
    wire \uu2.vbuf_w_addr_user.un459_ci_0_cascade_ ;
    wire \uu2.o_adder_vbuf_w_addr_user_8_cascade_ ;
    wire \INVuu2.w_addr_user_7C_net ;
    wire \uu2.un437_ci_3 ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \uu2.un2_w_addr_user_4_cascade_ ;
    wire \uu2.un2_w_addr_user_5 ;
    wire \uu2.un448_ci_5_cascade_ ;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \uu2.un415_ci ;
    wire \INVuu2.w_addr_user_5C_net ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire \uu2.mem0.w_addr_4 ;
    wire \uu2.mem0.g0_8_0_cascade_ ;
    wire \uu2.mem0.w_data_ns_1_1_0_3_cascade_ ;
    wire \uu2.Z_decfrac106 ;
    wire \uu2.mem0.w_data_ns_1_0_0_1_3 ;
    wire \uu2.g0_1_0_0_1_cascade_ ;
    wire \uu2.g0_1_0_0 ;
    wire \INVuu2.w_addr_displaying_5_rep1C_net ;
    wire \uu2.g0_1_a5_0_0 ;
    wire \uu2.g0_1_a5_1_0 ;
    wire \uu2.g1_1 ;
    wire \INVuu2.w_addr_displaying_2_rep1C_net ;
    wire \uu2.w_addr_displaying_8_repZ0Z1 ;
    wire \uu2.g1_0_1_cascade_ ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_50_cascade_ ;
    wire \uu2.g1_0_1 ;
    wire \uu2.mem0.g0_0 ;
    wire \uu2.w_addr_displaying_7_repZ0Z1 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_ ;
    wire \uu2.mem0.g1 ;
    wire \uu2.N_10 ;
    wire \uu2.mem0.g1_1_1 ;
    wire \INVuu2.w_addr_displaying_0_rep1C_net ;
    wire \uu2.w_addr_displaying_0_repZ0Z1 ;
    wire \uu2.mem0.N_10_0 ;
    wire \uu2.w_addr_displaying_4_rep1_3_cascade_ ;
    wire \uu2.w_addr_displaying_1_repZ0Z1 ;
    wire \uu2.w_addr_displaying_fastZ0Z_2 ;
    wire \uu2.mem0.un1_segment4_0_i_i_1 ;
    wire \INVuu2.w_addr_displaying_3_rep1C_net ;
    wire \uu2.mem0.un1_segment4_0_i_i_a5_0_0 ;
    wire \Lab_UT.didpuu0.didpsones.q13_0_cascade_ ;
    wire \uu2.g0_3Z0Z_0 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire bfn_7_14_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire \INVuu2.w_addr_user_0C_net ;
    wire \uu2.w_addr_user_2Z0Z_1_cascade_ ;
    wire \uu2.w_addr_userZ2Z_1_cascade_ ;
    wire \uu2.w_addr_user_RNIT1MGDZ0Z_4 ;
    wire \uu2.w_addr_user_1_0 ;
    wire \Lab_UT.dictrluu0.dek.det_NZ0Z_5_cascade_ ;
    wire \uu2.mem0.N_1476_0_0_0 ;
    wire \Lab_UT.dspStr.cnt11_1 ;
    wire \uu2.w_m5_i_a3Z0Z_2 ;
    wire \Lab_UT.dictrluu0.dek.det_NZ0Z_4 ;
    wire \uu2.un1_w_user_lf_0_0Z0Z_0_cascade_ ;
    wire \uu2.un1_w_user_lf_2 ;
    wire \uu2.un2_w_addr_user ;
    wire \uu2.un1_w_user_lf_2_cascade_ ;
    wire \uu2.un27_N_6_mux_0 ;
    wire CONSTANT_ONE_NET;
    wire \uu2.w_addr_user_RNILDNK6Z0Z_4_cascade_ ;
    wire \uu2.un27_w_addr_user_i ;
    wire \uu2.un1_w_user_lf_5_a0Z0Z_5_cascade_ ;
    wire \uu2.un1_w_user_lf_5_aZ0Z0 ;
    wire Lab_UT_dspStr_cnt_1_rep1;
    wire Lab_UT_dspStr_un36_dOut;
    wire Lab_UT_dspStr_un36_dOut_cascade_;
    wire \uu2.un27_N_6_mux_cascade_ ;
    wire \uu2.un27_w_addr_user_iZ0Z_1 ;
    wire Lab_UT_dspStr_cnt_3_rep1;
    wire Lab_UT_dspStr_cnt_2_rep1;
    wire L3_tx_data_0;
    wire L3_tx_data_0_cascade_;
    wire \uu2.un1_w_user_crZ0Z_1 ;
    wire \uu2.w_addr_displaying_RNIQKOV8Z0Z_8_cascade_ ;
    wire L3_tx_data_rdy;
    wire \uu2.un21_w_addr_displaying_i_cascade_ ;
    wire \INVuu2.w_addr_displaying_fast_6C_net ;
    wire \uu2.mem0.g0_i_a11_1_0 ;
    wire \uu2.w_addr_displaying_4_repZ0Z1 ;
    wire \uu2.mem0.g3_0_cascade_ ;
    wire \uu2.w_addr_displaying_3_repZ0Z1 ;
    wire \uu2.mem0.un1_segment4_0_i_i_0_0 ;
    wire \uu2.mem0.g0_i_a11_3_1 ;
    wire \uu2.mem0.g0_i_a11_7_1_cascade_ ;
    wire \uu2.mem0.g0_i_5_1 ;
    wire \INVuu2.w_addr_displaying_fast_0C_net ;
    wire \uu2.w_addr_displaying_fastZ0Z_0 ;
    wire \uu2.w_addr_displaying_6_repZ0Z1 ;
    wire \uu2.w_addr_displaying_5_repZ0Z1 ;
    wire \uu2.mem0.bitmap_pmux_1_1_i_a5_1_0 ;
    wire \uu2.mem0.g1_1_0_cascade_ ;
    wire \uu2.Z_decfrac106_5 ;
    wire \uu2.mem0.g0_2_0 ;
    wire \uu2.mem0.bitmap_pmux_1_1_i_a5_2_3_1_0 ;
    wire \uu2.w_addr_displaying_2_repZ0Z1 ;
    wire \uu2.Z_decfrac105_7_2 ;
    wire \uu2.w_addr_displaying_fastZ0Z_1 ;
    wire \INVuu2.w_addr_displaying_fast_1C_net ;
    wire \uu2.w_addr_displaying_fastZ0Z_4 ;
    wire \uu2.mem0.Z_decfrac105_7_3_2 ;
    wire \uu2.w_addr_displaying_4_8_cascade_ ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \uu2.un15_w_data_displaying ;
    wire \uu2.un15_w_data_displaying_cascade_ ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \uu2.w_addr_displaying_fastZ0Z_7 ;
    wire \INVuu2.w_addr_displaying_8C_net ;
    wire \uu2.un448_ci_5 ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire bfn_8_12_0_;
    wire \Lab_UT.didpuu0.didpsones.un1_q_cry_0 ;
    wire \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_2 ;
    wire \Lab_UT.didpuu0.didpsones.un1_q_cry_1 ;
    wire \Lab_UT.didpuu0.didpsones.un1_q_cry_2 ;
    wire \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_3_cascade_ ;
    wire \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_0 ;
    wire \Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_1 ;
    wire \Lab_UT.didpuu0.didpsones.q13_0 ;
    wire rst;
    wire \buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0 ;
    wire bfn_8_13_0_;
    wire \buart.Z_tx.bitcount_RNO_0Z0Z_1 ;
    wire \buart.Z_tx.un1_bitcount_cry_0 ;
    wire \buart.Z_tx.bitcount_RNO_0Z0Z_2 ;
    wire \buart.Z_tx.un1_bitcount_cry_1 ;
    wire uu2_un3_r_clk_en_0;
    wire \buart.Z_tx.un1_bitcount_cry_2 ;
    wire \buart.Z_tx.bitcount_RNIM5O32Z0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire buart__tx_uart_busy_0_cascade_;
    wire \buart.Z_tx.bitcount_RNIL4O32Z0Z_1 ;
    wire \buart.Z_tx.ser_clk ;
    wire buart__tx_uart_busy_0;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.un1_bitcount_axb_3 ;
    wire \Lab_UT.dspStr.cnt11_0_i ;
    wire \Lab_UT.dspStr.cntZ0Z_0 ;
    wire bfn_9_5_0_;
    wire \Lab_UT.dspStr.un1_cnt_3_cry_0 ;
    wire \Lab_UT.dspStr.un1_cnt_3_cry_1 ;
    wire \Lab_UT.dspStr.un1_cnt_3_cry_2 ;
    wire Lab_UT_dspStr_cnt_1;
    wire buart__rx_bitcount_3;
    wire buart__rx_bitcount_2;
    wire N_87;
    wire \Lab_UT.rx_data_rdy ;
    wire buart__rx_bitcount_0;
    wire \resetGen.un3_reset_count_i_a3Z0Z_4 ;
    wire Lab_UT_L3_tx_data_0_6;
    wire Lab_UT_dspStr_cnt_2;
    wire Lab_UT_dspStr_cnt_3;
    wire \Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9EZ0 ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.un4_w_user_data_rdyZ0Z_0 ;
    wire \uu2.mem0.w_addr_0 ;
    wire Lab_UT_L3_tx_data_0_5_cascade_;
    wire Lab_UT_L3_tx_data_0_2_6;
    wire \uu2.un1_w_user_crZ0Z_4 ;
    wire Lab_UT_L3_tx_data_0_2_1;
    wire Lab_UT_L3_tx_data_2_3;
    wire \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87EZ0 ;
    wire L3_tx_data_2;
    wire \Lab_UT.dspStr.cnt_fastZ0Z_1 ;
    wire \Lab_UT.dspStr.cnt_fastZ0Z_3 ;
    wire Lab_UT_L3_tx_data_0_4;
    wire \Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8EZ0 ;
    wire \Lab_UT.dspStr.cnt_fastZ0Z_2 ;
    wire Lab_UT_rx_data_0;
    wire Lab_UT_rx_data_1;
    wire Lab_UT_rx_data_2;
    wire Lab_UT_rx_data_3;
    wire Lab_UT_rx_data_6;
    wire \uu2.w_addr_displaying_fastZ0Z_6 ;
    wire \uu2.mem0.N_13_0 ;
    wire \uu2.w_addr_displayingZ0Z_3 ;
    wire \uu2.w_addr_displaying_4_3 ;
    wire Lab_UT_rx_data_7;
    wire Lab_UT_rx_data_5;
    wire Lab_UT_rx_data_4;
    wire \uu2.un1_w_user_lf_5_a0Z0Z_4 ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.un437_ci ;
    wire bu_rx_data_rdy;
    wire \Lab_UT.Lab3U00.bu_rx_data_rdy_0 ;
    wire \Lab_UT.sec_clkD ;
    wire \Lab_UT.didpuu0.clkSecStrbZ0 ;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \uu2.w_addr_displaying_fastZ0Z_3 ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \uu2.w_addr_displaying_4_fast_3 ;
    wire \uu2.mem0.g0_i_a11_2_0 ;
    wire \uu2.un15_w_data_displaying_5 ;
    wire \uu2.w_addr_displayingZ0Z_4 ;
    wire \uu2.w_addr_displaying_fastZ0Z_5 ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.un21_w_addr_displaying_i ;
    wire \uu2.w_addr_displaying_4_fast_8 ;
    wire \uu2.w_addr_displaying_fastZ0Z_8 ;
    wire \INVuu2.w_addr_displaying_fast_5C_net ;
    wire resetGen_rst_iso_g;
    wire \resetGen.un3_reset_count_i_a3Z0Z_5 ;
    wire bu_rx_data_0;
    wire bu_rx_data_1;
    wire bu_rx_data_7;
    wire bu_rx_data_6;
    wire bu_rx_data_5;
    wire bu_rx_data_4;
    wire bu_rx_data_3;
    wire bu_rx_data_2;
    wire clk_g;
    wire \buart.Z_rx.N_57_i ;
    wire Lab_UT_di_Sones_0;
    wire led_c_0;
    wire Lab_UT_dicRun;
    wire Lab_UT_l_oneSecPluse;
    wire led_c_4;
    wire Lab_UT_di_Sones_2;
    wire led_c_2;
    wire Lab_UT_di_Sones_3;
    wire led_c_3;
    wire \Lab_UT.dicSelectLEDdisp ;
    wire Lab_UT_di_Sones_1;
    wire led_c_1;
    wire _gnd_net_;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(latticehx1k_pll_inst_PLLOUTCORE_i),
            .REFERENCECLK(N__5054),
            .RESETB(N__8894),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__5510,N__5471,N__5495,N__5453,N__5423,N__5608,N__5639,N__5675,N__5579}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__5282,N__7898,N__5360,N__5252,N__7949,N__5237,N__5264,N__5273,N__11135}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,N__7316,dangling_wire_29,N__7355,dangling_wire_30,N__7667,dangling_wire_31,N__5243,dangling_wire_32,N__7724,dangling_wire_33,N__7634,dangling_wire_34,N__5375,dangling_wire_35,N__7646}),
            .RCLKE(N__5828),
            .RCLK(N__13421),
            .RE(N__5827),
            .WCLKE(N__7588),
            .WCLK(N__13420),
            .WE(N__7592));
    IO_PAD led_obuf_4_iopad (
            .OE(N__13611),
            .DIN(N__13610),
            .DOUT(N__13609),
            .PACKAGEPIN(led[4]));
    defparam led_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_4_preio (
            .PADOEN(N__13611),
            .PADOUT(N__13610),
            .PADIN(N__13609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13076),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__13602),
            .DIN(N__13601),
            .DOUT(N__13600),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__13602),
            .PADOUT(N__13601),
            .PADIN(N__13600),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_1_iopad (
            .OE(N__13593),
            .DIN(N__13592),
            .DOUT(N__13591),
            .PACKAGEPIN(led[1]));
    defparam led_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_1_preio (
            .PADOEN(N__13593),
            .PADOUT(N__13592),
            .PADIN(N__13591),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12818),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__13584),
            .DIN(N__13583),
            .DOUT(N__13582),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__13584),
            .PADOUT(N__13583),
            .PADIN(N__13582),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7187),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__13575),
            .DIN(N__13574),
            .DOUT(N__13573),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__13575),
            .PADOUT(N__13574),
            .PADIN(N__13573),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_2_iopad (
            .OE(N__13566),
            .DIN(N__13565),
            .DOUT(N__13564),
            .PACKAGEPIN(led[2]));
    defparam led_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_2_preio (
            .PADOEN(N__13566),
            .PADOUT(N__13565),
            .PADIN(N__13564),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13010),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_3_iopad (
            .OE(N__13557),
            .DIN(N__13556),
            .DOUT(N__13555),
            .PACKAGEPIN(led[3]));
    defparam led_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_3_preio (
            .PADOEN(N__13557),
            .PADOUT(N__13556),
            .PADIN(N__13555),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12932),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuf_0_iopad (
            .OE(N__13548),
            .DIN(N__13547),
            .DOUT(N__13546),
            .PACKAGEPIN(led[0]));
    defparam led_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO led_obuf_0_preio (
            .PADOEN(N__13548),
            .PADOUT(N__13547),
            .PADIN(N__13546),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13178),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__13539),
            .DIN(N__13538),
            .DOUT(N__13537),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__13539),
            .PADOUT(N__13538),
            .PADIN(N__13537),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__13415),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__13530),
            .DIN(N__13529),
            .DOUT(N__13528),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__13530),
            .PADOUT(N__13529),
            .PADIN(N__13528),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__3253 (
            .O(N__13511),
            .I(N__13507));
    InMux I__3252 (
            .O(N__13510),
            .I(N__13503));
    LocalMux I__3251 (
            .O(N__13507),
            .I(N__13500));
    InMux I__3250 (
            .O(N__13506),
            .I(N__13497));
    LocalMux I__3249 (
            .O(N__13503),
            .I(N__13492));
    Span4Mux_v I__3248 (
            .O(N__13500),
            .I(N__13492));
    LocalMux I__3247 (
            .O(N__13497),
            .I(bu_rx_data_4));
    Odrv4 I__3246 (
            .O(N__13492),
            .I(bu_rx_data_4));
    InMux I__3245 (
            .O(N__13487),
            .I(N__13483));
    InMux I__3244 (
            .O(N__13486),
            .I(N__13480));
    LocalMux I__3243 (
            .O(N__13483),
            .I(N__13474));
    LocalMux I__3242 (
            .O(N__13480),
            .I(N__13474));
    InMux I__3241 (
            .O(N__13479),
            .I(N__13471));
    Span4Mux_v I__3240 (
            .O(N__13474),
            .I(N__13468));
    LocalMux I__3239 (
            .O(N__13471),
            .I(bu_rx_data_3));
    Odrv4 I__3238 (
            .O(N__13468),
            .I(bu_rx_data_3));
    InMux I__3237 (
            .O(N__13463),
            .I(N__13459));
    InMux I__3236 (
            .O(N__13462),
            .I(N__13456));
    LocalMux I__3235 (
            .O(N__13459),
            .I(N__13453));
    LocalMux I__3234 (
            .O(N__13456),
            .I(N__13449));
    Span4Mux_v I__3233 (
            .O(N__13453),
            .I(N__13446));
    InMux I__3232 (
            .O(N__13452),
            .I(N__13443));
    Span4Mux_v I__3231 (
            .O(N__13449),
            .I(N__13438));
    Span4Mux_h I__3230 (
            .O(N__13446),
            .I(N__13438));
    LocalMux I__3229 (
            .O(N__13443),
            .I(bu_rx_data_2));
    Odrv4 I__3228 (
            .O(N__13438),
            .I(bu_rx_data_2));
    ClkMux I__3227 (
            .O(N__13433),
            .I(N__13265));
    ClkMux I__3226 (
            .O(N__13432),
            .I(N__13265));
    ClkMux I__3225 (
            .O(N__13431),
            .I(N__13265));
    ClkMux I__3224 (
            .O(N__13430),
            .I(N__13265));
    ClkMux I__3223 (
            .O(N__13429),
            .I(N__13265));
    ClkMux I__3222 (
            .O(N__13428),
            .I(N__13265));
    ClkMux I__3221 (
            .O(N__13427),
            .I(N__13265));
    ClkMux I__3220 (
            .O(N__13426),
            .I(N__13265));
    ClkMux I__3219 (
            .O(N__13425),
            .I(N__13265));
    ClkMux I__3218 (
            .O(N__13424),
            .I(N__13265));
    ClkMux I__3217 (
            .O(N__13423),
            .I(N__13265));
    ClkMux I__3216 (
            .O(N__13422),
            .I(N__13265));
    ClkMux I__3215 (
            .O(N__13421),
            .I(N__13265));
    ClkMux I__3214 (
            .O(N__13420),
            .I(N__13265));
    ClkMux I__3213 (
            .O(N__13419),
            .I(N__13265));
    ClkMux I__3212 (
            .O(N__13418),
            .I(N__13265));
    ClkMux I__3211 (
            .O(N__13417),
            .I(N__13265));
    ClkMux I__3210 (
            .O(N__13416),
            .I(N__13265));
    ClkMux I__3209 (
            .O(N__13415),
            .I(N__13265));
    ClkMux I__3208 (
            .O(N__13414),
            .I(N__13265));
    ClkMux I__3207 (
            .O(N__13413),
            .I(N__13265));
    ClkMux I__3206 (
            .O(N__13412),
            .I(N__13265));
    ClkMux I__3205 (
            .O(N__13411),
            .I(N__13265));
    ClkMux I__3204 (
            .O(N__13410),
            .I(N__13265));
    ClkMux I__3203 (
            .O(N__13409),
            .I(N__13265));
    ClkMux I__3202 (
            .O(N__13408),
            .I(N__13265));
    ClkMux I__3201 (
            .O(N__13407),
            .I(N__13265));
    ClkMux I__3200 (
            .O(N__13406),
            .I(N__13265));
    ClkMux I__3199 (
            .O(N__13405),
            .I(N__13265));
    ClkMux I__3198 (
            .O(N__13404),
            .I(N__13265));
    ClkMux I__3197 (
            .O(N__13403),
            .I(N__13265));
    ClkMux I__3196 (
            .O(N__13402),
            .I(N__13265));
    ClkMux I__3195 (
            .O(N__13401),
            .I(N__13265));
    ClkMux I__3194 (
            .O(N__13400),
            .I(N__13265));
    ClkMux I__3193 (
            .O(N__13399),
            .I(N__13265));
    ClkMux I__3192 (
            .O(N__13398),
            .I(N__13265));
    ClkMux I__3191 (
            .O(N__13397),
            .I(N__13265));
    ClkMux I__3190 (
            .O(N__13396),
            .I(N__13265));
    ClkMux I__3189 (
            .O(N__13395),
            .I(N__13265));
    ClkMux I__3188 (
            .O(N__13394),
            .I(N__13265));
    ClkMux I__3187 (
            .O(N__13393),
            .I(N__13265));
    ClkMux I__3186 (
            .O(N__13392),
            .I(N__13265));
    ClkMux I__3185 (
            .O(N__13391),
            .I(N__13265));
    ClkMux I__3184 (
            .O(N__13390),
            .I(N__13265));
    ClkMux I__3183 (
            .O(N__13389),
            .I(N__13265));
    ClkMux I__3182 (
            .O(N__13388),
            .I(N__13265));
    ClkMux I__3181 (
            .O(N__13387),
            .I(N__13265));
    ClkMux I__3180 (
            .O(N__13386),
            .I(N__13265));
    ClkMux I__3179 (
            .O(N__13385),
            .I(N__13265));
    ClkMux I__3178 (
            .O(N__13384),
            .I(N__13265));
    ClkMux I__3177 (
            .O(N__13383),
            .I(N__13265));
    ClkMux I__3176 (
            .O(N__13382),
            .I(N__13265));
    ClkMux I__3175 (
            .O(N__13381),
            .I(N__13265));
    ClkMux I__3174 (
            .O(N__13380),
            .I(N__13265));
    ClkMux I__3173 (
            .O(N__13379),
            .I(N__13265));
    ClkMux I__3172 (
            .O(N__13378),
            .I(N__13265));
    GlobalMux I__3171 (
            .O(N__13265),
            .I(N__13262));
    gio2CtrlBuf I__3170 (
            .O(N__13262),
            .I(clk_g));
    CEMux I__3169 (
            .O(N__13259),
            .I(N__13256));
    LocalMux I__3168 (
            .O(N__13256),
            .I(N__13252));
    CEMux I__3167 (
            .O(N__13255),
            .I(N__13249));
    Span4Mux_v I__3166 (
            .O(N__13252),
            .I(N__13246));
    LocalMux I__3165 (
            .O(N__13249),
            .I(N__13243));
    Span4Mux_s2_h I__3164 (
            .O(N__13246),
            .I(N__13240));
    Span4Mux_v I__3163 (
            .O(N__13243),
            .I(N__13237));
    Odrv4 I__3162 (
            .O(N__13240),
            .I(\buart.Z_rx.N_57_i ));
    Odrv4 I__3161 (
            .O(N__13237),
            .I(\buart.Z_rx.N_57_i ));
    InMux I__3160 (
            .O(N__13232),
            .I(N__13229));
    LocalMux I__3159 (
            .O(N__13229),
            .I(N__13220));
    InMux I__3158 (
            .O(N__13228),
            .I(N__13211));
    InMux I__3157 (
            .O(N__13227),
            .I(N__13211));
    InMux I__3156 (
            .O(N__13226),
            .I(N__13211));
    InMux I__3155 (
            .O(N__13225),
            .I(N__13211));
    InMux I__3154 (
            .O(N__13224),
            .I(N__13205));
    InMux I__3153 (
            .O(N__13223),
            .I(N__13202));
    Span4Mux_v I__3152 (
            .O(N__13220),
            .I(N__13199));
    LocalMux I__3151 (
            .O(N__13211),
            .I(N__13196));
    InMux I__3150 (
            .O(N__13210),
            .I(N__13189));
    InMux I__3149 (
            .O(N__13209),
            .I(N__13189));
    InMux I__3148 (
            .O(N__13208),
            .I(N__13189));
    LocalMux I__3147 (
            .O(N__13205),
            .I(Lab_UT_di_Sones_0));
    LocalMux I__3146 (
            .O(N__13202),
            .I(Lab_UT_di_Sones_0));
    Odrv4 I__3145 (
            .O(N__13199),
            .I(Lab_UT_di_Sones_0));
    Odrv12 I__3144 (
            .O(N__13196),
            .I(Lab_UT_di_Sones_0));
    LocalMux I__3143 (
            .O(N__13189),
            .I(Lab_UT_di_Sones_0));
    IoInMux I__3142 (
            .O(N__13178),
            .I(N__13175));
    LocalMux I__3141 (
            .O(N__13175),
            .I(N__13172));
    Odrv12 I__3140 (
            .O(N__13172),
            .I(led_c_0));
    InMux I__3139 (
            .O(N__13169),
            .I(N__13165));
    InMux I__3138 (
            .O(N__13168),
            .I(N__13162));
    LocalMux I__3137 (
            .O(N__13165),
            .I(N__13155));
    LocalMux I__3136 (
            .O(N__13162),
            .I(N__13155));
    InMux I__3135 (
            .O(N__13161),
            .I(N__13150));
    InMux I__3134 (
            .O(N__13160),
            .I(N__13150));
    Odrv12 I__3133 (
            .O(N__13155),
            .I(Lab_UT_dicRun));
    LocalMux I__3132 (
            .O(N__13150),
            .I(Lab_UT_dicRun));
    CascadeMux I__3131 (
            .O(N__13145),
            .I(N__13141));
    InMux I__3130 (
            .O(N__13144),
            .I(N__13137));
    InMux I__3129 (
            .O(N__13141),
            .I(N__13131));
    InMux I__3128 (
            .O(N__13140),
            .I(N__13131));
    LocalMux I__3127 (
            .O(N__13137),
            .I(N__13128));
    InMux I__3126 (
            .O(N__13136),
            .I(N__13125));
    LocalMux I__3125 (
            .O(N__13131),
            .I(N__13122));
    Span4Mux_v I__3124 (
            .O(N__13128),
            .I(N__13118));
    LocalMux I__3123 (
            .O(N__13125),
            .I(N__13114));
    Span4Mux_h I__3122 (
            .O(N__13122),
            .I(N__13111));
    InMux I__3121 (
            .O(N__13121),
            .I(N__13108));
    Span4Mux_v I__3120 (
            .O(N__13118),
            .I(N__13104));
    InMux I__3119 (
            .O(N__13117),
            .I(N__13101));
    Span4Mux_v I__3118 (
            .O(N__13114),
            .I(N__13094));
    Span4Mux_v I__3117 (
            .O(N__13111),
            .I(N__13094));
    LocalMux I__3116 (
            .O(N__13108),
            .I(N__13094));
    InMux I__3115 (
            .O(N__13107),
            .I(N__13091));
    Sp12to4 I__3114 (
            .O(N__13104),
            .I(N__13086));
    LocalMux I__3113 (
            .O(N__13101),
            .I(N__13086));
    Span4Mux_h I__3112 (
            .O(N__13094),
            .I(N__13083));
    LocalMux I__3111 (
            .O(N__13091),
            .I(Lab_UT_l_oneSecPluse));
    Odrv12 I__3110 (
            .O(N__13086),
            .I(Lab_UT_l_oneSecPluse));
    Odrv4 I__3109 (
            .O(N__13083),
            .I(Lab_UT_l_oneSecPluse));
    IoInMux I__3108 (
            .O(N__13076),
            .I(N__13073));
    LocalMux I__3107 (
            .O(N__13073),
            .I(N__13070));
    Odrv4 I__3106 (
            .O(N__13070),
            .I(led_c_4));
    InMux I__3105 (
            .O(N__13067),
            .I(N__13062));
    CascadeMux I__3104 (
            .O(N__13066),
            .I(N__13059));
    CascadeMux I__3103 (
            .O(N__13065),
            .I(N__13056));
    LocalMux I__3102 (
            .O(N__13062),
            .I(N__13051));
    InMux I__3101 (
            .O(N__13059),
            .I(N__13044));
    InMux I__3100 (
            .O(N__13056),
            .I(N__13044));
    InMux I__3099 (
            .O(N__13055),
            .I(N__13044));
    InMux I__3098 (
            .O(N__13054),
            .I(N__13041));
    Span4Mux_v I__3097 (
            .O(N__13051),
            .I(N__13033));
    LocalMux I__3096 (
            .O(N__13044),
            .I(N__13033));
    LocalMux I__3095 (
            .O(N__13041),
            .I(N__13033));
    InMux I__3094 (
            .O(N__13040),
            .I(N__13027));
    Span4Mux_h I__3093 (
            .O(N__13033),
            .I(N__13024));
    InMux I__3092 (
            .O(N__13032),
            .I(N__13017));
    InMux I__3091 (
            .O(N__13031),
            .I(N__13017));
    InMux I__3090 (
            .O(N__13030),
            .I(N__13017));
    LocalMux I__3089 (
            .O(N__13027),
            .I(Lab_UT_di_Sones_2));
    Odrv4 I__3088 (
            .O(N__13024),
            .I(Lab_UT_di_Sones_2));
    LocalMux I__3087 (
            .O(N__13017),
            .I(Lab_UT_di_Sones_2));
    IoInMux I__3086 (
            .O(N__13010),
            .I(N__13007));
    LocalMux I__3085 (
            .O(N__13007),
            .I(N__13004));
    Odrv4 I__3084 (
            .O(N__13004),
            .I(led_c_2));
    InMux I__3083 (
            .O(N__13001),
            .I(N__12995));
    CascadeMux I__3082 (
            .O(N__13000),
            .I(N__12992));
    CascadeMux I__3081 (
            .O(N__12999),
            .I(N__12988));
    CascadeMux I__3080 (
            .O(N__12998),
            .I(N__12985));
    LocalMux I__3079 (
            .O(N__12995),
            .I(N__12980));
    InMux I__3078 (
            .O(N__12992),
            .I(N__12976));
    InMux I__3077 (
            .O(N__12991),
            .I(N__12967));
    InMux I__3076 (
            .O(N__12988),
            .I(N__12967));
    InMux I__3075 (
            .O(N__12985),
            .I(N__12967));
    InMux I__3074 (
            .O(N__12984),
            .I(N__12967));
    CascadeMux I__3073 (
            .O(N__12983),
            .I(N__12963));
    Span4Mux_h I__3072 (
            .O(N__12980),
            .I(N__12959));
    InMux I__3071 (
            .O(N__12979),
            .I(N__12956));
    LocalMux I__3070 (
            .O(N__12976),
            .I(N__12953));
    LocalMux I__3069 (
            .O(N__12967),
            .I(N__12950));
    InMux I__3068 (
            .O(N__12966),
            .I(N__12943));
    InMux I__3067 (
            .O(N__12963),
            .I(N__12943));
    InMux I__3066 (
            .O(N__12962),
            .I(N__12943));
    Odrv4 I__3065 (
            .O(N__12959),
            .I(Lab_UT_di_Sones_3));
    LocalMux I__3064 (
            .O(N__12956),
            .I(Lab_UT_di_Sones_3));
    Odrv4 I__3063 (
            .O(N__12953),
            .I(Lab_UT_di_Sones_3));
    Odrv12 I__3062 (
            .O(N__12950),
            .I(Lab_UT_di_Sones_3));
    LocalMux I__3061 (
            .O(N__12943),
            .I(Lab_UT_di_Sones_3));
    IoInMux I__3060 (
            .O(N__12932),
            .I(N__12929));
    LocalMux I__3059 (
            .O(N__12929),
            .I(N__12926));
    Odrv4 I__3058 (
            .O(N__12926),
            .I(led_c_3));
    InMux I__3057 (
            .O(N__12923),
            .I(N__12920));
    LocalMux I__3056 (
            .O(N__12920),
            .I(N__12916));
    InMux I__3055 (
            .O(N__12919),
            .I(N__12911));
    Span4Mux_v I__3054 (
            .O(N__12916),
            .I(N__12908));
    InMux I__3053 (
            .O(N__12915),
            .I(N__12903));
    InMux I__3052 (
            .O(N__12914),
            .I(N__12903));
    LocalMux I__3051 (
            .O(N__12911),
            .I(N__12900));
    Sp12to4 I__3050 (
            .O(N__12908),
            .I(N__12895));
    LocalMux I__3049 (
            .O(N__12903),
            .I(N__12895));
    Span4Mux_v I__3048 (
            .O(N__12900),
            .I(N__12892));
    Span12Mux_s4_h I__3047 (
            .O(N__12895),
            .I(N__12889));
    Span4Mux_v I__3046 (
            .O(N__12892),
            .I(N__12886));
    Odrv12 I__3045 (
            .O(N__12889),
            .I(\Lab_UT.dicSelectLEDdisp ));
    Odrv4 I__3044 (
            .O(N__12886),
            .I(\Lab_UT.dicSelectLEDdisp ));
    InMux I__3043 (
            .O(N__12881),
            .I(N__12877));
    InMux I__3042 (
            .O(N__12880),
            .I(N__12868));
    LocalMux I__3041 (
            .O(N__12877),
            .I(N__12864));
    CascadeMux I__3040 (
            .O(N__12876),
            .I(N__12861));
    CascadeMux I__3039 (
            .O(N__12875),
            .I(N__12857));
    InMux I__3038 (
            .O(N__12874),
            .I(N__12848));
    InMux I__3037 (
            .O(N__12873),
            .I(N__12848));
    InMux I__3036 (
            .O(N__12872),
            .I(N__12848));
    InMux I__3035 (
            .O(N__12871),
            .I(N__12848));
    LocalMux I__3034 (
            .O(N__12868),
            .I(N__12845));
    InMux I__3033 (
            .O(N__12867),
            .I(N__12842));
    Span4Mux_s3_h I__3032 (
            .O(N__12864),
            .I(N__12839));
    InMux I__3031 (
            .O(N__12861),
            .I(N__12832));
    InMux I__3030 (
            .O(N__12860),
            .I(N__12832));
    InMux I__3029 (
            .O(N__12857),
            .I(N__12832));
    LocalMux I__3028 (
            .O(N__12848),
            .I(N__12829));
    Odrv12 I__3027 (
            .O(N__12845),
            .I(Lab_UT_di_Sones_1));
    LocalMux I__3026 (
            .O(N__12842),
            .I(Lab_UT_di_Sones_1));
    Odrv4 I__3025 (
            .O(N__12839),
            .I(Lab_UT_di_Sones_1));
    LocalMux I__3024 (
            .O(N__12832),
            .I(Lab_UT_di_Sones_1));
    Odrv12 I__3023 (
            .O(N__12829),
            .I(Lab_UT_di_Sones_1));
    IoInMux I__3022 (
            .O(N__12818),
            .I(N__12815));
    LocalMux I__3021 (
            .O(N__12815),
            .I(N__12812));
    Odrv4 I__3020 (
            .O(N__12812),
            .I(led_c_1));
    CascadeMux I__3019 (
            .O(N__12809),
            .I(N__12805));
    CascadeMux I__3018 (
            .O(N__12808),
            .I(N__12799));
    InMux I__3017 (
            .O(N__12805),
            .I(N__12793));
    InMux I__3016 (
            .O(N__12804),
            .I(N__12788));
    InMux I__3015 (
            .O(N__12803),
            .I(N__12784));
    InMux I__3014 (
            .O(N__12802),
            .I(N__12777));
    InMux I__3013 (
            .O(N__12799),
            .I(N__12777));
    InMux I__3012 (
            .O(N__12798),
            .I(N__12777));
    CascadeMux I__3011 (
            .O(N__12797),
            .I(N__12774));
    CascadeMux I__3010 (
            .O(N__12796),
            .I(N__12770));
    LocalMux I__3009 (
            .O(N__12793),
            .I(N__12766));
    InMux I__3008 (
            .O(N__12792),
            .I(N__12763));
    InMux I__3007 (
            .O(N__12791),
            .I(N__12760));
    LocalMux I__3006 (
            .O(N__12788),
            .I(N__12756));
    InMux I__3005 (
            .O(N__12787),
            .I(N__12753));
    LocalMux I__3004 (
            .O(N__12784),
            .I(N__12748));
    LocalMux I__3003 (
            .O(N__12777),
            .I(N__12748));
    InMux I__3002 (
            .O(N__12774),
            .I(N__12739));
    InMux I__3001 (
            .O(N__12773),
            .I(N__12739));
    InMux I__3000 (
            .O(N__12770),
            .I(N__12739));
    InMux I__2999 (
            .O(N__12769),
            .I(N__12739));
    Span4Mux_h I__2998 (
            .O(N__12766),
            .I(N__12732));
    LocalMux I__2997 (
            .O(N__12763),
            .I(N__12732));
    LocalMux I__2996 (
            .O(N__12760),
            .I(N__12732));
    InMux I__2995 (
            .O(N__12759),
            .I(N__12729));
    Span12Mux_s8_v I__2994 (
            .O(N__12756),
            .I(N__12726));
    LocalMux I__2993 (
            .O(N__12753),
            .I(N__12719));
    Span4Mux_h I__2992 (
            .O(N__12748),
            .I(N__12719));
    LocalMux I__2991 (
            .O(N__12739),
            .I(N__12719));
    Odrv4 I__2990 (
            .O(N__12732),
            .I(\uu2.un15_w_data_displaying_5 ));
    LocalMux I__2989 (
            .O(N__12729),
            .I(\uu2.un15_w_data_displaying_5 ));
    Odrv12 I__2988 (
            .O(N__12726),
            .I(\uu2.un15_w_data_displaying_5 ));
    Odrv4 I__2987 (
            .O(N__12719),
            .I(\uu2.un15_w_data_displaying_5 ));
    InMux I__2986 (
            .O(N__12710),
            .I(N__12707));
    LocalMux I__2985 (
            .O(N__12707),
            .I(N__12702));
    InMux I__2984 (
            .O(N__12706),
            .I(N__12699));
    CascadeMux I__2983 (
            .O(N__12705),
            .I(N__12695));
    Span4Mux_v I__2982 (
            .O(N__12702),
            .I(N__12687));
    LocalMux I__2981 (
            .O(N__12699),
            .I(N__12687));
    CascadeMux I__2980 (
            .O(N__12698),
            .I(N__12678));
    InMux I__2979 (
            .O(N__12695),
            .I(N__12672));
    InMux I__2978 (
            .O(N__12694),
            .I(N__12669));
    InMux I__2977 (
            .O(N__12693),
            .I(N__12664));
    InMux I__2976 (
            .O(N__12692),
            .I(N__12664));
    Span4Mux_h I__2975 (
            .O(N__12687),
            .I(N__12661));
    InMux I__2974 (
            .O(N__12686),
            .I(N__12658));
    InMux I__2973 (
            .O(N__12685),
            .I(N__12651));
    InMux I__2972 (
            .O(N__12684),
            .I(N__12651));
    InMux I__2971 (
            .O(N__12683),
            .I(N__12651));
    InMux I__2970 (
            .O(N__12682),
            .I(N__12644));
    InMux I__2969 (
            .O(N__12681),
            .I(N__12644));
    InMux I__2968 (
            .O(N__12678),
            .I(N__12644));
    InMux I__2967 (
            .O(N__12677),
            .I(N__12637));
    InMux I__2966 (
            .O(N__12676),
            .I(N__12637));
    InMux I__2965 (
            .O(N__12675),
            .I(N__12637));
    LocalMux I__2964 (
            .O(N__12672),
            .I(N__12634));
    LocalMux I__2963 (
            .O(N__12669),
            .I(N__12629));
    LocalMux I__2962 (
            .O(N__12664),
            .I(N__12629));
    Odrv4 I__2961 (
            .O(N__12661),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2960 (
            .O(N__12658),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2959 (
            .O(N__12651),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2958 (
            .O(N__12644),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2957 (
            .O(N__12637),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv12 I__2956 (
            .O(N__12634),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2955 (
            .O(N__12629),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    InMux I__2954 (
            .O(N__12614),
            .I(N__12610));
    InMux I__2953 (
            .O(N__12613),
            .I(N__12607));
    LocalMux I__2952 (
            .O(N__12610),
            .I(\uu2.w_addr_displaying_fastZ0Z_5 ));
    LocalMux I__2951 (
            .O(N__12607),
            .I(\uu2.w_addr_displaying_fastZ0Z_5 ));
    CascadeMux I__2950 (
            .O(N__12602),
            .I(N__12595));
    CascadeMux I__2949 (
            .O(N__12601),
            .I(N__12592));
    CascadeMux I__2948 (
            .O(N__12600),
            .I(N__12587));
    InMux I__2947 (
            .O(N__12599),
            .I(N__12581));
    InMux I__2946 (
            .O(N__12598),
            .I(N__12576));
    InMux I__2945 (
            .O(N__12595),
            .I(N__12576));
    InMux I__2944 (
            .O(N__12592),
            .I(N__12567));
    InMux I__2943 (
            .O(N__12591),
            .I(N__12567));
    InMux I__2942 (
            .O(N__12590),
            .I(N__12567));
    InMux I__2941 (
            .O(N__12587),
            .I(N__12567));
    InMux I__2940 (
            .O(N__12586),
            .I(N__12564));
    CascadeMux I__2939 (
            .O(N__12585),
            .I(N__12558));
    InMux I__2938 (
            .O(N__12584),
            .I(N__12555));
    LocalMux I__2937 (
            .O(N__12581),
            .I(N__12550));
    LocalMux I__2936 (
            .O(N__12576),
            .I(N__12550));
    LocalMux I__2935 (
            .O(N__12567),
            .I(N__12547));
    LocalMux I__2934 (
            .O(N__12564),
            .I(N__12544));
    InMux I__2933 (
            .O(N__12563),
            .I(N__12541));
    InMux I__2932 (
            .O(N__12562),
            .I(N__12538));
    InMux I__2931 (
            .O(N__12561),
            .I(N__12533));
    InMux I__2930 (
            .O(N__12558),
            .I(N__12533));
    LocalMux I__2929 (
            .O(N__12555),
            .I(N__12530));
    Span4Mux_v I__2928 (
            .O(N__12550),
            .I(N__12525));
    Span4Mux_v I__2927 (
            .O(N__12547),
            .I(N__12525));
    Span4Mux_h I__2926 (
            .O(N__12544),
            .I(N__12522));
    LocalMux I__2925 (
            .O(N__12541),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2924 (
            .O(N__12538),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2923 (
            .O(N__12533),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv12 I__2922 (
            .O(N__12530),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__2921 (
            .O(N__12525),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__2920 (
            .O(N__12522),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    CascadeMux I__2919 (
            .O(N__12509),
            .I(N__12505));
    CascadeMux I__2918 (
            .O(N__12508),
            .I(N__12490));
    InMux I__2917 (
            .O(N__12505),
            .I(N__12476));
    InMux I__2916 (
            .O(N__12504),
            .I(N__12476));
    InMux I__2915 (
            .O(N__12503),
            .I(N__12476));
    InMux I__2914 (
            .O(N__12502),
            .I(N__12476));
    InMux I__2913 (
            .O(N__12501),
            .I(N__12469));
    InMux I__2912 (
            .O(N__12500),
            .I(N__12469));
    InMux I__2911 (
            .O(N__12499),
            .I(N__12469));
    InMux I__2910 (
            .O(N__12498),
            .I(N__12457));
    InMux I__2909 (
            .O(N__12497),
            .I(N__12457));
    InMux I__2908 (
            .O(N__12496),
            .I(N__12450));
    InMux I__2907 (
            .O(N__12495),
            .I(N__12450));
    InMux I__2906 (
            .O(N__12494),
            .I(N__12450));
    InMux I__2905 (
            .O(N__12493),
            .I(N__12447));
    InMux I__2904 (
            .O(N__12490),
            .I(N__12442));
    InMux I__2903 (
            .O(N__12489),
            .I(N__12442));
    InMux I__2902 (
            .O(N__12488),
            .I(N__12433));
    InMux I__2901 (
            .O(N__12487),
            .I(N__12433));
    InMux I__2900 (
            .O(N__12486),
            .I(N__12433));
    InMux I__2899 (
            .O(N__12485),
            .I(N__12433));
    LocalMux I__2898 (
            .O(N__12476),
            .I(N__12428));
    LocalMux I__2897 (
            .O(N__12469),
            .I(N__12428));
    InMux I__2896 (
            .O(N__12468),
            .I(N__12423));
    InMux I__2895 (
            .O(N__12467),
            .I(N__12423));
    InMux I__2894 (
            .O(N__12466),
            .I(N__12420));
    InMux I__2893 (
            .O(N__12465),
            .I(N__12417));
    InMux I__2892 (
            .O(N__12464),
            .I(N__12410));
    InMux I__2891 (
            .O(N__12463),
            .I(N__12410));
    InMux I__2890 (
            .O(N__12462),
            .I(N__12410));
    LocalMux I__2889 (
            .O(N__12457),
            .I(N__12407));
    LocalMux I__2888 (
            .O(N__12450),
            .I(N__12404));
    LocalMux I__2887 (
            .O(N__12447),
            .I(N__12401));
    LocalMux I__2886 (
            .O(N__12442),
            .I(N__12394));
    LocalMux I__2885 (
            .O(N__12433),
            .I(N__12394));
    Span4Mux_h I__2884 (
            .O(N__12428),
            .I(N__12394));
    LocalMux I__2883 (
            .O(N__12423),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__2882 (
            .O(N__12420),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__2881 (
            .O(N__12417),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__2880 (
            .O(N__12410),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__2879 (
            .O(N__12407),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__2878 (
            .O(N__12404),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__2877 (
            .O(N__12401),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__2876 (
            .O(N__12394),
            .I(\uu2.un21_w_addr_displaying_i ));
    InMux I__2875 (
            .O(N__12377),
            .I(N__12374));
    LocalMux I__2874 (
            .O(N__12374),
            .I(\uu2.w_addr_displaying_4_fast_8 ));
    CascadeMux I__2873 (
            .O(N__12371),
            .I(N__12367));
    InMux I__2872 (
            .O(N__12370),
            .I(N__12362));
    InMux I__2871 (
            .O(N__12367),
            .I(N__12362));
    LocalMux I__2870 (
            .O(N__12362),
            .I(N__12359));
    Span4Mux_h I__2869 (
            .O(N__12359),
            .I(N__12352));
    CascadeMux I__2868 (
            .O(N__12358),
            .I(N__12349));
    CascadeMux I__2867 (
            .O(N__12357),
            .I(N__12346));
    InMux I__2866 (
            .O(N__12356),
            .I(N__12343));
    InMux I__2865 (
            .O(N__12355),
            .I(N__12340));
    Span4Mux_s3_h I__2864 (
            .O(N__12352),
            .I(N__12337));
    InMux I__2863 (
            .O(N__12349),
            .I(N__12332));
    InMux I__2862 (
            .O(N__12346),
            .I(N__12332));
    LocalMux I__2861 (
            .O(N__12343),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    LocalMux I__2860 (
            .O(N__12340),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    Odrv4 I__2859 (
            .O(N__12337),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    LocalMux I__2858 (
            .O(N__12332),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    InMux I__2857 (
            .O(N__12323),
            .I(N__12318));
    SRMux I__2856 (
            .O(N__12322),
            .I(N__12313));
    InMux I__2855 (
            .O(N__12321),
            .I(N__12313));
    LocalMux I__2854 (
            .O(N__12318),
            .I(N__12295));
    LocalMux I__2853 (
            .O(N__12313),
            .I(N__12292));
    SRMux I__2852 (
            .O(N__12312),
            .I(N__12224));
    SRMux I__2851 (
            .O(N__12311),
            .I(N__12224));
    SRMux I__2850 (
            .O(N__12310),
            .I(N__12224));
    SRMux I__2849 (
            .O(N__12309),
            .I(N__12224));
    SRMux I__2848 (
            .O(N__12308),
            .I(N__12224));
    SRMux I__2847 (
            .O(N__12307),
            .I(N__12224));
    SRMux I__2846 (
            .O(N__12306),
            .I(N__12224));
    SRMux I__2845 (
            .O(N__12305),
            .I(N__12224));
    SRMux I__2844 (
            .O(N__12304),
            .I(N__12224));
    SRMux I__2843 (
            .O(N__12303),
            .I(N__12224));
    SRMux I__2842 (
            .O(N__12302),
            .I(N__12224));
    SRMux I__2841 (
            .O(N__12301),
            .I(N__12224));
    SRMux I__2840 (
            .O(N__12300),
            .I(N__12224));
    SRMux I__2839 (
            .O(N__12299),
            .I(N__12224));
    SRMux I__2838 (
            .O(N__12298),
            .I(N__12224));
    Glb2LocalMux I__2837 (
            .O(N__12295),
            .I(N__12224));
    Glb2LocalMux I__2836 (
            .O(N__12292),
            .I(N__12224));
    SRMux I__2835 (
            .O(N__12291),
            .I(N__12224));
    SRMux I__2834 (
            .O(N__12290),
            .I(N__12224));
    SRMux I__2833 (
            .O(N__12289),
            .I(N__12224));
    SRMux I__2832 (
            .O(N__12288),
            .I(N__12224));
    SRMux I__2831 (
            .O(N__12287),
            .I(N__12224));
    SRMux I__2830 (
            .O(N__12286),
            .I(N__12224));
    SRMux I__2829 (
            .O(N__12285),
            .I(N__12224));
    SRMux I__2828 (
            .O(N__12284),
            .I(N__12224));
    SRMux I__2827 (
            .O(N__12283),
            .I(N__12224));
    SRMux I__2826 (
            .O(N__12282),
            .I(N__12224));
    SRMux I__2825 (
            .O(N__12281),
            .I(N__12224));
    GlobalMux I__2824 (
            .O(N__12224),
            .I(N__12221));
    gio2CtrlBuf I__2823 (
            .O(N__12221),
            .I(resetGen_rst_iso_g));
    InMux I__2822 (
            .O(N__12218),
            .I(N__12215));
    LocalMux I__2821 (
            .O(N__12215),
            .I(N__12212));
    Span4Mux_h I__2820 (
            .O(N__12212),
            .I(N__12209));
    Odrv4 I__2819 (
            .O(N__12209),
            .I(\resetGen.un3_reset_count_i_a3Z0Z_5 ));
    InMux I__2818 (
            .O(N__12206),
            .I(N__12203));
    LocalMux I__2817 (
            .O(N__12203),
            .I(N__12199));
    InMux I__2816 (
            .O(N__12202),
            .I(N__12196));
    Odrv4 I__2815 (
            .O(N__12199),
            .I(bu_rx_data_0));
    LocalMux I__2814 (
            .O(N__12196),
            .I(bu_rx_data_0));
    InMux I__2813 (
            .O(N__12191),
            .I(N__12188));
    LocalMux I__2812 (
            .O(N__12188),
            .I(N__12183));
    InMux I__2811 (
            .O(N__12187),
            .I(N__12178));
    InMux I__2810 (
            .O(N__12186),
            .I(N__12178));
    Odrv4 I__2809 (
            .O(N__12183),
            .I(bu_rx_data_1));
    LocalMux I__2808 (
            .O(N__12178),
            .I(bu_rx_data_1));
    InMux I__2807 (
            .O(N__12173),
            .I(N__12169));
    CascadeMux I__2806 (
            .O(N__12172),
            .I(N__12165));
    LocalMux I__2805 (
            .O(N__12169),
            .I(N__12162));
    InMux I__2804 (
            .O(N__12168),
            .I(N__12159));
    InMux I__2803 (
            .O(N__12165),
            .I(N__12156));
    Span4Mux_s3_h I__2802 (
            .O(N__12162),
            .I(N__12151));
    LocalMux I__2801 (
            .O(N__12159),
            .I(N__12151));
    LocalMux I__2800 (
            .O(N__12156),
            .I(N__12148));
    Span4Mux_v I__2799 (
            .O(N__12151),
            .I(N__12145));
    Span4Mux_v I__2798 (
            .O(N__12148),
            .I(N__12142));
    Odrv4 I__2797 (
            .O(N__12145),
            .I(bu_rx_data_7));
    Odrv4 I__2796 (
            .O(N__12142),
            .I(bu_rx_data_7));
    InMux I__2795 (
            .O(N__12137),
            .I(N__12133));
    CascadeMux I__2794 (
            .O(N__12136),
            .I(N__12129));
    LocalMux I__2793 (
            .O(N__12133),
            .I(N__12126));
    InMux I__2792 (
            .O(N__12132),
            .I(N__12121));
    InMux I__2791 (
            .O(N__12129),
            .I(N__12121));
    Odrv4 I__2790 (
            .O(N__12126),
            .I(bu_rx_data_6));
    LocalMux I__2789 (
            .O(N__12121),
            .I(bu_rx_data_6));
    InMux I__2788 (
            .O(N__12116),
            .I(N__12113));
    LocalMux I__2787 (
            .O(N__12113),
            .I(N__12108));
    InMux I__2786 (
            .O(N__12112),
            .I(N__12103));
    InMux I__2785 (
            .O(N__12111),
            .I(N__12103));
    Odrv12 I__2784 (
            .O(N__12108),
            .I(bu_rx_data_5));
    LocalMux I__2783 (
            .O(N__12103),
            .I(bu_rx_data_5));
    InMux I__2782 (
            .O(N__12098),
            .I(N__12094));
    InMux I__2781 (
            .O(N__12097),
            .I(N__12091));
    LocalMux I__2780 (
            .O(N__12094),
            .I(\uu2.w_addr_displaying_fastZ0Z_6 ));
    LocalMux I__2779 (
            .O(N__12091),
            .I(\uu2.w_addr_displaying_fastZ0Z_6 ));
    InMux I__2778 (
            .O(N__12086),
            .I(N__12083));
    LocalMux I__2777 (
            .O(N__12083),
            .I(\uu2.mem0.N_13_0 ));
    InMux I__2776 (
            .O(N__12080),
            .I(N__12074));
    InMux I__2775 (
            .O(N__12079),
            .I(N__12069));
    CascadeMux I__2774 (
            .O(N__12078),
            .I(N__12066));
    InMux I__2773 (
            .O(N__12077),
            .I(N__12060));
    LocalMux I__2772 (
            .O(N__12074),
            .I(N__12056));
    InMux I__2771 (
            .O(N__12073),
            .I(N__12051));
    InMux I__2770 (
            .O(N__12072),
            .I(N__12051));
    LocalMux I__2769 (
            .O(N__12069),
            .I(N__12046));
    InMux I__2768 (
            .O(N__12066),
            .I(N__12043));
    InMux I__2767 (
            .O(N__12065),
            .I(N__12038));
    InMux I__2766 (
            .O(N__12064),
            .I(N__12038));
    InMux I__2765 (
            .O(N__12063),
            .I(N__12035));
    LocalMux I__2764 (
            .O(N__12060),
            .I(N__12032));
    InMux I__2763 (
            .O(N__12059),
            .I(N__12029));
    Span4Mux_v I__2762 (
            .O(N__12056),
            .I(N__12024));
    LocalMux I__2761 (
            .O(N__12051),
            .I(N__12024));
    InMux I__2760 (
            .O(N__12050),
            .I(N__12019));
    InMux I__2759 (
            .O(N__12049),
            .I(N__12019));
    Span4Mux_h I__2758 (
            .O(N__12046),
            .I(N__12012));
    LocalMux I__2757 (
            .O(N__12043),
            .I(N__12012));
    LocalMux I__2756 (
            .O(N__12038),
            .I(N__12012));
    LocalMux I__2755 (
            .O(N__12035),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2754 (
            .O(N__12032),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2753 (
            .O(N__12029),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2752 (
            .O(N__12024),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2751 (
            .O(N__12019),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2750 (
            .O(N__12012),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    InMux I__2749 (
            .O(N__11999),
            .I(N__11996));
    LocalMux I__2748 (
            .O(N__11996),
            .I(N__11993));
    Span4Mux_v I__2747 (
            .O(N__11993),
            .I(N__11990));
    Span4Mux_h I__2746 (
            .O(N__11990),
            .I(N__11987));
    Odrv4 I__2745 (
            .O(N__11987),
            .I(\uu2.w_addr_displaying_4_3 ));
    InMux I__2744 (
            .O(N__11984),
            .I(N__11979));
    InMux I__2743 (
            .O(N__11983),
            .I(N__11974));
    InMux I__2742 (
            .O(N__11982),
            .I(N__11974));
    LocalMux I__2741 (
            .O(N__11979),
            .I(N__11971));
    LocalMux I__2740 (
            .O(N__11974),
            .I(N__11968));
    Span4Mux_h I__2739 (
            .O(N__11971),
            .I(N__11963));
    Span4Mux_h I__2738 (
            .O(N__11968),
            .I(N__11960));
    InMux I__2737 (
            .O(N__11967),
            .I(N__11957));
    InMux I__2736 (
            .O(N__11966),
            .I(N__11954));
    Odrv4 I__2735 (
            .O(N__11963),
            .I(Lab_UT_rx_data_7));
    Odrv4 I__2734 (
            .O(N__11960),
            .I(Lab_UT_rx_data_7));
    LocalMux I__2733 (
            .O(N__11957),
            .I(Lab_UT_rx_data_7));
    LocalMux I__2732 (
            .O(N__11954),
            .I(Lab_UT_rx_data_7));
    CascadeMux I__2731 (
            .O(N__11945),
            .I(N__11941));
    InMux I__2730 (
            .O(N__11944),
            .I(N__11938));
    InMux I__2729 (
            .O(N__11941),
            .I(N__11935));
    LocalMux I__2728 (
            .O(N__11938),
            .I(N__11931));
    LocalMux I__2727 (
            .O(N__11935),
            .I(N__11928));
    InMux I__2726 (
            .O(N__11934),
            .I(N__11925));
    Span4Mux_h I__2725 (
            .O(N__11931),
            .I(N__11919));
    Span4Mux_h I__2724 (
            .O(N__11928),
            .I(N__11919));
    LocalMux I__2723 (
            .O(N__11925),
            .I(N__11916));
    InMux I__2722 (
            .O(N__11924),
            .I(N__11913));
    Odrv4 I__2721 (
            .O(N__11919),
            .I(Lab_UT_rx_data_5));
    Odrv4 I__2720 (
            .O(N__11916),
            .I(Lab_UT_rx_data_5));
    LocalMux I__2719 (
            .O(N__11913),
            .I(Lab_UT_rx_data_5));
    InMux I__2718 (
            .O(N__11906),
            .I(N__11900));
    InMux I__2717 (
            .O(N__11905),
            .I(N__11900));
    LocalMux I__2716 (
            .O(N__11900),
            .I(N__11895));
    InMux I__2715 (
            .O(N__11899),
            .I(N__11892));
    InMux I__2714 (
            .O(N__11898),
            .I(N__11889));
    Odrv4 I__2713 (
            .O(N__11895),
            .I(Lab_UT_rx_data_4));
    LocalMux I__2712 (
            .O(N__11892),
            .I(Lab_UT_rx_data_4));
    LocalMux I__2711 (
            .O(N__11889),
            .I(Lab_UT_rx_data_4));
    InMux I__2710 (
            .O(N__11882),
            .I(N__11879));
    LocalMux I__2709 (
            .O(N__11879),
            .I(N__11876));
    Odrv4 I__2708 (
            .O(N__11876),
            .I(\uu2.un1_w_user_lf_5_a0Z0Z_4 ));
    InMux I__2707 (
            .O(N__11873),
            .I(N__11869));
    InMux I__2706 (
            .O(N__11872),
            .I(N__11866));
    LocalMux I__2705 (
            .O(N__11869),
            .I(N__11860));
    LocalMux I__2704 (
            .O(N__11866),
            .I(N__11857));
    InMux I__2703 (
            .O(N__11865),
            .I(N__11852));
    InMux I__2702 (
            .O(N__11864),
            .I(N__11852));
    CascadeMux I__2701 (
            .O(N__11863),
            .I(N__11849));
    Span4Mux_v I__2700 (
            .O(N__11860),
            .I(N__11840));
    Span4Mux_v I__2699 (
            .O(N__11857),
            .I(N__11840));
    LocalMux I__2698 (
            .O(N__11852),
            .I(N__11840));
    InMux I__2697 (
            .O(N__11849),
            .I(N__11835));
    InMux I__2696 (
            .O(N__11848),
            .I(N__11835));
    InMux I__2695 (
            .O(N__11847),
            .I(N__11832));
    Odrv4 I__2694 (
            .O(N__11840),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2693 (
            .O(N__11835),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2692 (
            .O(N__11832),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    CascadeMux I__2691 (
            .O(N__11825),
            .I(N__11822));
    InMux I__2690 (
            .O(N__11822),
            .I(N__11819));
    LocalMux I__2689 (
            .O(N__11819),
            .I(N__11814));
    InMux I__2688 (
            .O(N__11818),
            .I(N__11811));
    InMux I__2687 (
            .O(N__11817),
            .I(N__11808));
    Span4Mux_h I__2686 (
            .O(N__11814),
            .I(N__11803));
    LocalMux I__2685 (
            .O(N__11811),
            .I(N__11803));
    LocalMux I__2684 (
            .O(N__11808),
            .I(N__11800));
    Odrv4 I__2683 (
            .O(N__11803),
            .I(\uu2.un437_ci ));
    Odrv4 I__2682 (
            .O(N__11800),
            .I(\uu2.un437_ci ));
    InMux I__2681 (
            .O(N__11795),
            .I(N__11791));
    InMux I__2680 (
            .O(N__11794),
            .I(N__11788));
    LocalMux I__2679 (
            .O(N__11791),
            .I(N__11785));
    LocalMux I__2678 (
            .O(N__11788),
            .I(N__11782));
    Span4Mux_v I__2677 (
            .O(N__11785),
            .I(N__11778));
    Span4Mux_h I__2676 (
            .O(N__11782),
            .I(N__11775));
    InMux I__2675 (
            .O(N__11781),
            .I(N__11772));
    Odrv4 I__2674 (
            .O(N__11778),
            .I(bu_rx_data_rdy));
    Odrv4 I__2673 (
            .O(N__11775),
            .I(bu_rx_data_rdy));
    LocalMux I__2672 (
            .O(N__11772),
            .I(bu_rx_data_rdy));
    CEMux I__2671 (
            .O(N__11765),
            .I(N__11762));
    LocalMux I__2670 (
            .O(N__11762),
            .I(N__11759));
    Odrv12 I__2669 (
            .O(N__11759),
            .I(\Lab_UT.Lab3U00.bu_rx_data_rdy_0 ));
    CascadeMux I__2668 (
            .O(N__11756),
            .I(N__11752));
    InMux I__2667 (
            .O(N__11755),
            .I(N__11749));
    InMux I__2666 (
            .O(N__11752),
            .I(N__11746));
    LocalMux I__2665 (
            .O(N__11749),
            .I(N__11743));
    LocalMux I__2664 (
            .O(N__11746),
            .I(N__11740));
    Span4Mux_v I__2663 (
            .O(N__11743),
            .I(N__11735));
    Span4Mux_h I__2662 (
            .O(N__11740),
            .I(N__11735));
    Odrv4 I__2661 (
            .O(N__11735),
            .I(\Lab_UT.sec_clkD ));
    InMux I__2660 (
            .O(N__11732),
            .I(N__11726));
    InMux I__2659 (
            .O(N__11731),
            .I(N__11721));
    InMux I__2658 (
            .O(N__11730),
            .I(N__11721));
    CascadeMux I__2657 (
            .O(N__11729),
            .I(N__11716));
    LocalMux I__2656 (
            .O(N__11726),
            .I(N__11711));
    LocalMux I__2655 (
            .O(N__11721),
            .I(N__11711));
    InMux I__2654 (
            .O(N__11720),
            .I(N__11704));
    InMux I__2653 (
            .O(N__11719),
            .I(N__11704));
    InMux I__2652 (
            .O(N__11716),
            .I(N__11704));
    Span4Mux_h I__2651 (
            .O(N__11711),
            .I(N__11699));
    LocalMux I__2650 (
            .O(N__11704),
            .I(N__11699));
    Odrv4 I__2649 (
            .O(N__11699),
            .I(\Lab_UT.didpuu0.clkSecStrbZ0 ));
    InMux I__2648 (
            .O(N__11696),
            .I(N__11687));
    InMux I__2647 (
            .O(N__11695),
            .I(N__11687));
    InMux I__2646 (
            .O(N__11694),
            .I(N__11684));
    InMux I__2645 (
            .O(N__11693),
            .I(N__11678));
    InMux I__2644 (
            .O(N__11692),
            .I(N__11678));
    LocalMux I__2643 (
            .O(N__11687),
            .I(N__11671));
    LocalMux I__2642 (
            .O(N__11684),
            .I(N__11668));
    InMux I__2641 (
            .O(N__11683),
            .I(N__11665));
    LocalMux I__2640 (
            .O(N__11678),
            .I(N__11662));
    InMux I__2639 (
            .O(N__11677),
            .I(N__11653));
    InMux I__2638 (
            .O(N__11676),
            .I(N__11653));
    InMux I__2637 (
            .O(N__11675),
            .I(N__11653));
    InMux I__2636 (
            .O(N__11674),
            .I(N__11653));
    Span4Mux_s3_h I__2635 (
            .O(N__11671),
            .I(N__11646));
    Span4Mux_v I__2634 (
            .O(N__11668),
            .I(N__11646));
    LocalMux I__2633 (
            .O(N__11665),
            .I(N__11646));
    Odrv4 I__2632 (
            .O(N__11662),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__2631 (
            .O(N__11653),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__2630 (
            .O(N__11646),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    CascadeMux I__2629 (
            .O(N__11639),
            .I(N__11634));
    CascadeMux I__2628 (
            .O(N__11638),
            .I(N__11630));
    CascadeMux I__2627 (
            .O(N__11637),
            .I(N__11624));
    InMux I__2626 (
            .O(N__11634),
            .I(N__11621));
    InMux I__2625 (
            .O(N__11633),
            .I(N__11618));
    InMux I__2624 (
            .O(N__11630),
            .I(N__11609));
    InMux I__2623 (
            .O(N__11629),
            .I(N__11609));
    InMux I__2622 (
            .O(N__11628),
            .I(N__11609));
    InMux I__2621 (
            .O(N__11627),
            .I(N__11609));
    InMux I__2620 (
            .O(N__11624),
            .I(N__11606));
    LocalMux I__2619 (
            .O(N__11621),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__2618 (
            .O(N__11618),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__2617 (
            .O(N__11609),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__2616 (
            .O(N__11606),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    CascadeMux I__2615 (
            .O(N__11597),
            .I(N__11593));
    InMux I__2614 (
            .O(N__11596),
            .I(N__11587));
    InMux I__2613 (
            .O(N__11593),
            .I(N__11583));
    CascadeMux I__2612 (
            .O(N__11592),
            .I(N__11580));
    InMux I__2611 (
            .O(N__11591),
            .I(N__11575));
    InMux I__2610 (
            .O(N__11590),
            .I(N__11575));
    LocalMux I__2609 (
            .O(N__11587),
            .I(N__11572));
    InMux I__2608 (
            .O(N__11586),
            .I(N__11568));
    LocalMux I__2607 (
            .O(N__11583),
            .I(N__11565));
    InMux I__2606 (
            .O(N__11580),
            .I(N__11561));
    LocalMux I__2605 (
            .O(N__11575),
            .I(N__11558));
    Span4Mux_h I__2604 (
            .O(N__11572),
            .I(N__11555));
    InMux I__2603 (
            .O(N__11571),
            .I(N__11552));
    LocalMux I__2602 (
            .O(N__11568),
            .I(N__11547));
    Span4Mux_h I__2601 (
            .O(N__11565),
            .I(N__11547));
    InMux I__2600 (
            .O(N__11564),
            .I(N__11544));
    LocalMux I__2599 (
            .O(N__11561),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2598 (
            .O(N__11558),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2597 (
            .O(N__11555),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__2596 (
            .O(N__11552),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2595 (
            .O(N__11547),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__2594 (
            .O(N__11544),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    InMux I__2593 (
            .O(N__11531),
            .I(N__11528));
    LocalMux I__2592 (
            .O(N__11528),
            .I(N__11525));
    Odrv4 I__2591 (
            .O(N__11525),
            .I(\uu2.w_addr_displaying_4_fast_3 ));
    InMux I__2590 (
            .O(N__11522),
            .I(N__11519));
    LocalMux I__2589 (
            .O(N__11519),
            .I(N__11516));
    Odrv4 I__2588 (
            .O(N__11516),
            .I(\uu2.mem0.g0_i_a11_2_0 ));
    InMux I__2587 (
            .O(N__11513),
            .I(N__11510));
    LocalMux I__2586 (
            .O(N__11510),
            .I(N__11506));
    InMux I__2585 (
            .O(N__11509),
            .I(N__11503));
    Sp12to4 I__2584 (
            .O(N__11506),
            .I(N__11497));
    LocalMux I__2583 (
            .O(N__11503),
            .I(N__11497));
    InMux I__2582 (
            .O(N__11502),
            .I(N__11494));
    Odrv12 I__2581 (
            .O(N__11497),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8EZ0 ));
    LocalMux I__2580 (
            .O(N__11494),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8EZ0 ));
    CascadeMux I__2579 (
            .O(N__11489),
            .I(N__11484));
    CascadeMux I__2578 (
            .O(N__11488),
            .I(N__11480));
    CascadeMux I__2577 (
            .O(N__11487),
            .I(N__11477));
    InMux I__2576 (
            .O(N__11484),
            .I(N__11465));
    InMux I__2575 (
            .O(N__11483),
            .I(N__11465));
    InMux I__2574 (
            .O(N__11480),
            .I(N__11465));
    InMux I__2573 (
            .O(N__11477),
            .I(N__11465));
    InMux I__2572 (
            .O(N__11476),
            .I(N__11465));
    LocalMux I__2571 (
            .O(N__11465),
            .I(\Lab_UT.dspStr.cnt_fastZ0Z_2 ));
    InMux I__2570 (
            .O(N__11462),
            .I(N__11459));
    LocalMux I__2569 (
            .O(N__11459),
            .I(N__11452));
    CascadeMux I__2568 (
            .O(N__11458),
            .I(N__11449));
    InMux I__2567 (
            .O(N__11457),
            .I(N__11445));
    InMux I__2566 (
            .O(N__11456),
            .I(N__11440));
    InMux I__2565 (
            .O(N__11455),
            .I(N__11440));
    Span4Mux_h I__2564 (
            .O(N__11452),
            .I(N__11437));
    InMux I__2563 (
            .O(N__11449),
            .I(N__11432));
    InMux I__2562 (
            .O(N__11448),
            .I(N__11432));
    LocalMux I__2561 (
            .O(N__11445),
            .I(N__11427));
    LocalMux I__2560 (
            .O(N__11440),
            .I(N__11427));
    Odrv4 I__2559 (
            .O(N__11437),
            .I(Lab_UT_rx_data_0));
    LocalMux I__2558 (
            .O(N__11432),
            .I(Lab_UT_rx_data_0));
    Odrv4 I__2557 (
            .O(N__11427),
            .I(Lab_UT_rx_data_0));
    CascadeMux I__2556 (
            .O(N__11420),
            .I(N__11417));
    InMux I__2555 (
            .O(N__11417),
            .I(N__11413));
    InMux I__2554 (
            .O(N__11416),
            .I(N__11410));
    LocalMux I__2553 (
            .O(N__11413),
            .I(N__11405));
    LocalMux I__2552 (
            .O(N__11410),
            .I(N__11402));
    InMux I__2551 (
            .O(N__11409),
            .I(N__11399));
    InMux I__2550 (
            .O(N__11408),
            .I(N__11396));
    Odrv4 I__2549 (
            .O(N__11405),
            .I(Lab_UT_rx_data_1));
    Odrv12 I__2548 (
            .O(N__11402),
            .I(Lab_UT_rx_data_1));
    LocalMux I__2547 (
            .O(N__11399),
            .I(Lab_UT_rx_data_1));
    LocalMux I__2546 (
            .O(N__11396),
            .I(Lab_UT_rx_data_1));
    InMux I__2545 (
            .O(N__11387),
            .I(N__11383));
    InMux I__2544 (
            .O(N__11386),
            .I(N__11379));
    LocalMux I__2543 (
            .O(N__11383),
            .I(N__11375));
    InMux I__2542 (
            .O(N__11382),
            .I(N__11372));
    LocalMux I__2541 (
            .O(N__11379),
            .I(N__11369));
    InMux I__2540 (
            .O(N__11378),
            .I(N__11366));
    Odrv4 I__2539 (
            .O(N__11375),
            .I(Lab_UT_rx_data_2));
    LocalMux I__2538 (
            .O(N__11372),
            .I(Lab_UT_rx_data_2));
    Odrv4 I__2537 (
            .O(N__11369),
            .I(Lab_UT_rx_data_2));
    LocalMux I__2536 (
            .O(N__11366),
            .I(Lab_UT_rx_data_2));
    InMux I__2535 (
            .O(N__11357),
            .I(N__11351));
    InMux I__2534 (
            .O(N__11356),
            .I(N__11344));
    InMux I__2533 (
            .O(N__11355),
            .I(N__11344));
    InMux I__2532 (
            .O(N__11354),
            .I(N__11344));
    LocalMux I__2531 (
            .O(N__11351),
            .I(N__11338));
    LocalMux I__2530 (
            .O(N__11344),
            .I(N__11338));
    InMux I__2529 (
            .O(N__11343),
            .I(N__11335));
    Odrv4 I__2528 (
            .O(N__11338),
            .I(Lab_UT_rx_data_3));
    LocalMux I__2527 (
            .O(N__11335),
            .I(Lab_UT_rx_data_3));
    InMux I__2526 (
            .O(N__11330),
            .I(N__11324));
    InMux I__2525 (
            .O(N__11329),
            .I(N__11324));
    LocalMux I__2524 (
            .O(N__11324),
            .I(N__11320));
    CascadeMux I__2523 (
            .O(N__11323),
            .I(N__11317));
    Span4Mux_h I__2522 (
            .O(N__11320),
            .I(N__11314));
    InMux I__2521 (
            .O(N__11317),
            .I(N__11311));
    Odrv4 I__2520 (
            .O(N__11314),
            .I(Lab_UT_rx_data_6));
    LocalMux I__2519 (
            .O(N__11311),
            .I(Lab_UT_rx_data_6));
    InMux I__2518 (
            .O(N__11306),
            .I(N__11303));
    LocalMux I__2517 (
            .O(N__11303),
            .I(N__11300));
    Span4Mux_v I__2516 (
            .O(N__11300),
            .I(N__11295));
    InMux I__2515 (
            .O(N__11299),
            .I(N__11290));
    InMux I__2514 (
            .O(N__11298),
            .I(N__11290));
    Odrv4 I__2513 (
            .O(N__11295),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9EZ0 ));
    LocalMux I__2512 (
            .O(N__11290),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9EZ0 ));
    InMux I__2511 (
            .O(N__11285),
            .I(N__11281));
    InMux I__2510 (
            .O(N__11284),
            .I(N__11273));
    LocalMux I__2509 (
            .O(N__11281),
            .I(N__11270));
    InMux I__2508 (
            .O(N__11280),
            .I(N__11259));
    InMux I__2507 (
            .O(N__11279),
            .I(N__11259));
    InMux I__2506 (
            .O(N__11278),
            .I(N__11259));
    InMux I__2505 (
            .O(N__11277),
            .I(N__11259));
    InMux I__2504 (
            .O(N__11276),
            .I(N__11259));
    LocalMux I__2503 (
            .O(N__11273),
            .I(\uu2.w_addr_userZ0Z_0 ));
    Odrv4 I__2502 (
            .O(N__11270),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__2501 (
            .O(N__11259),
            .I(\uu2.w_addr_userZ0Z_0 ));
    InMux I__2500 (
            .O(N__11252),
            .I(N__11237));
    InMux I__2499 (
            .O(N__11251),
            .I(N__11237));
    InMux I__2498 (
            .O(N__11250),
            .I(N__11224));
    InMux I__2497 (
            .O(N__11249),
            .I(N__11224));
    InMux I__2496 (
            .O(N__11248),
            .I(N__11224));
    InMux I__2495 (
            .O(N__11247),
            .I(N__11224));
    InMux I__2494 (
            .O(N__11246),
            .I(N__11224));
    InMux I__2493 (
            .O(N__11245),
            .I(N__11224));
    CascadeMux I__2492 (
            .O(N__11244),
            .I(N__11221));
    InMux I__2491 (
            .O(N__11243),
            .I(N__11214));
    InMux I__2490 (
            .O(N__11242),
            .I(N__11210));
    LocalMux I__2489 (
            .O(N__11237),
            .I(N__11205));
    LocalMux I__2488 (
            .O(N__11224),
            .I(N__11205));
    InMux I__2487 (
            .O(N__11221),
            .I(N__11202));
    InMux I__2486 (
            .O(N__11220),
            .I(N__11198));
    InMux I__2485 (
            .O(N__11219),
            .I(N__11193));
    InMux I__2484 (
            .O(N__11218),
            .I(N__11193));
    InMux I__2483 (
            .O(N__11217),
            .I(N__11190));
    LocalMux I__2482 (
            .O(N__11214),
            .I(N__11187));
    InMux I__2481 (
            .O(N__11213),
            .I(N__11184));
    LocalMux I__2480 (
            .O(N__11210),
            .I(N__11180));
    Span4Mux_v I__2479 (
            .O(N__11205),
            .I(N__11175));
    LocalMux I__2478 (
            .O(N__11202),
            .I(N__11175));
    InMux I__2477 (
            .O(N__11201),
            .I(N__11172));
    LocalMux I__2476 (
            .O(N__11198),
            .I(N__11169));
    LocalMux I__2475 (
            .O(N__11193),
            .I(N__11166));
    LocalMux I__2474 (
            .O(N__11190),
            .I(N__11161));
    Span4Mux_h I__2473 (
            .O(N__11187),
            .I(N__11161));
    LocalMux I__2472 (
            .O(N__11184),
            .I(N__11158));
    InMux I__2471 (
            .O(N__11183),
            .I(N__11155));
    Span4Mux_h I__2470 (
            .O(N__11180),
            .I(N__11150));
    Span4Mux_h I__2469 (
            .O(N__11175),
            .I(N__11150));
    LocalMux I__2468 (
            .O(N__11172),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__2467 (
            .O(N__11169),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv12 I__2466 (
            .O(N__11166),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__2465 (
            .O(N__11161),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__2464 (
            .O(N__11158),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    LocalMux I__2463 (
            .O(N__11155),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__2462 (
            .O(N__11150),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    CascadeMux I__2461 (
            .O(N__11135),
            .I(N__11132));
    InMux I__2460 (
            .O(N__11132),
            .I(N__11129));
    LocalMux I__2459 (
            .O(N__11129),
            .I(N__11126));
    Span4Mux_h I__2458 (
            .O(N__11126),
            .I(N__11123));
    Span4Mux_h I__2457 (
            .O(N__11123),
            .I(N__11120));
    Odrv4 I__2456 (
            .O(N__11120),
            .I(\uu2.mem0.w_addr_0 ));
    CascadeMux I__2455 (
            .O(N__11117),
            .I(Lab_UT_L3_tx_data_0_5_cascade_));
    InMux I__2454 (
            .O(N__11114),
            .I(N__11110));
    InMux I__2453 (
            .O(N__11113),
            .I(N__11107));
    LocalMux I__2452 (
            .O(N__11110),
            .I(Lab_UT_L3_tx_data_0_2_6));
    LocalMux I__2451 (
            .O(N__11107),
            .I(Lab_UT_L3_tx_data_0_2_6));
    InMux I__2450 (
            .O(N__11102),
            .I(N__11096));
    InMux I__2449 (
            .O(N__11101),
            .I(N__11096));
    LocalMux I__2448 (
            .O(N__11096),
            .I(N__11092));
    InMux I__2447 (
            .O(N__11095),
            .I(N__11089));
    Span4Mux_h I__2446 (
            .O(N__11092),
            .I(N__11083));
    LocalMux I__2445 (
            .O(N__11089),
            .I(N__11080));
    InMux I__2444 (
            .O(N__11088),
            .I(N__11073));
    InMux I__2443 (
            .O(N__11087),
            .I(N__11073));
    InMux I__2442 (
            .O(N__11086),
            .I(N__11073));
    Odrv4 I__2441 (
            .O(N__11083),
            .I(\uu2.un1_w_user_crZ0Z_4 ));
    Odrv4 I__2440 (
            .O(N__11080),
            .I(\uu2.un1_w_user_crZ0Z_4 ));
    LocalMux I__2439 (
            .O(N__11073),
            .I(\uu2.un1_w_user_crZ0Z_4 ));
    InMux I__2438 (
            .O(N__11066),
            .I(N__11063));
    LocalMux I__2437 (
            .O(N__11063),
            .I(Lab_UT_L3_tx_data_0_2_1));
    InMux I__2436 (
            .O(N__11060),
            .I(N__11057));
    LocalMux I__2435 (
            .O(N__11057),
            .I(Lab_UT_L3_tx_data_2_3));
    InMux I__2434 (
            .O(N__11054),
            .I(N__11050));
    InMux I__2433 (
            .O(N__11053),
            .I(N__11047));
    LocalMux I__2432 (
            .O(N__11050),
            .I(N__11043));
    LocalMux I__2431 (
            .O(N__11047),
            .I(N__11040));
    InMux I__2430 (
            .O(N__11046),
            .I(N__11037));
    Odrv4 I__2429 (
            .O(N__11043),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87EZ0 ));
    Odrv4 I__2428 (
            .O(N__11040),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87EZ0 ));
    LocalMux I__2427 (
            .O(N__11037),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87EZ0 ));
    InMux I__2426 (
            .O(N__11030),
            .I(N__11027));
    LocalMux I__2425 (
            .O(N__11027),
            .I(N__11024));
    Span4Mux_h I__2424 (
            .O(N__11024),
            .I(N__11020));
    InMux I__2423 (
            .O(N__11023),
            .I(N__11017));
    Odrv4 I__2422 (
            .O(N__11020),
            .I(L3_tx_data_2));
    LocalMux I__2421 (
            .O(N__11017),
            .I(L3_tx_data_2));
    CascadeMux I__2420 (
            .O(N__11012),
            .I(N__11009));
    InMux I__2419 (
            .O(N__11009),
            .I(N__11002));
    InMux I__2418 (
            .O(N__11008),
            .I(N__10993));
    InMux I__2417 (
            .O(N__11007),
            .I(N__10993));
    InMux I__2416 (
            .O(N__11006),
            .I(N__10993));
    InMux I__2415 (
            .O(N__11005),
            .I(N__10993));
    LocalMux I__2414 (
            .O(N__11002),
            .I(\Lab_UT.dspStr.cnt_fastZ0Z_1 ));
    LocalMux I__2413 (
            .O(N__10993),
            .I(\Lab_UT.dspStr.cnt_fastZ0Z_1 ));
    CascadeMux I__2412 (
            .O(N__10988),
            .I(N__10981));
    InMux I__2411 (
            .O(N__10987),
            .I(N__10970));
    InMux I__2410 (
            .O(N__10986),
            .I(N__10970));
    InMux I__2409 (
            .O(N__10985),
            .I(N__10970));
    InMux I__2408 (
            .O(N__10984),
            .I(N__10970));
    InMux I__2407 (
            .O(N__10981),
            .I(N__10970));
    LocalMux I__2406 (
            .O(N__10970),
            .I(\Lab_UT.dspStr.cnt_fastZ0Z_3 ));
    InMux I__2405 (
            .O(N__10967),
            .I(N__10964));
    LocalMux I__2404 (
            .O(N__10964),
            .I(N__10960));
    InMux I__2403 (
            .O(N__10963),
            .I(N__10957));
    Odrv12 I__2402 (
            .O(N__10960),
            .I(Lab_UT_L3_tx_data_0_4));
    LocalMux I__2401 (
            .O(N__10957),
            .I(Lab_UT_L3_tx_data_0_4));
    InMux I__2400 (
            .O(N__10952),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_0 ));
    InMux I__2399 (
            .O(N__10949),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_1 ));
    InMux I__2398 (
            .O(N__10946),
            .I(\Lab_UT.dspStr.un1_cnt_3_cry_2 ));
    InMux I__2397 (
            .O(N__10943),
            .I(N__10937));
    InMux I__2396 (
            .O(N__10942),
            .I(N__10937));
    LocalMux I__2395 (
            .O(N__10937),
            .I(N__10932));
    InMux I__2394 (
            .O(N__10936),
            .I(N__10929));
    InMux I__2393 (
            .O(N__10935),
            .I(N__10926));
    Span4Mux_v I__2392 (
            .O(N__10932),
            .I(N__10921));
    LocalMux I__2391 (
            .O(N__10929),
            .I(N__10911));
    LocalMux I__2390 (
            .O(N__10926),
            .I(N__10911));
    InMux I__2389 (
            .O(N__10925),
            .I(N__10908));
    InMux I__2388 (
            .O(N__10924),
            .I(N__10905));
    Span4Mux_h I__2387 (
            .O(N__10921),
            .I(N__10902));
    InMux I__2386 (
            .O(N__10920),
            .I(N__10895));
    InMux I__2385 (
            .O(N__10919),
            .I(N__10895));
    InMux I__2384 (
            .O(N__10918),
            .I(N__10895));
    InMux I__2383 (
            .O(N__10917),
            .I(N__10890));
    InMux I__2382 (
            .O(N__10916),
            .I(N__10890));
    Span4Mux_h I__2381 (
            .O(N__10911),
            .I(N__10885));
    LocalMux I__2380 (
            .O(N__10908),
            .I(N__10885));
    LocalMux I__2379 (
            .O(N__10905),
            .I(Lab_UT_dspStr_cnt_1));
    Odrv4 I__2378 (
            .O(N__10902),
            .I(Lab_UT_dspStr_cnt_1));
    LocalMux I__2377 (
            .O(N__10895),
            .I(Lab_UT_dspStr_cnt_1));
    LocalMux I__2376 (
            .O(N__10890),
            .I(Lab_UT_dspStr_cnt_1));
    Odrv4 I__2375 (
            .O(N__10885),
            .I(Lab_UT_dspStr_cnt_1));
    InMux I__2374 (
            .O(N__10874),
            .I(N__10869));
    CascadeMux I__2373 (
            .O(N__10873),
            .I(N__10864));
    CascadeMux I__2372 (
            .O(N__10872),
            .I(N__10860));
    LocalMux I__2371 (
            .O(N__10869),
            .I(N__10856));
    InMux I__2370 (
            .O(N__10868),
            .I(N__10853));
    InMux I__2369 (
            .O(N__10867),
            .I(N__10850));
    InMux I__2368 (
            .O(N__10864),
            .I(N__10847));
    InMux I__2367 (
            .O(N__10863),
            .I(N__10840));
    InMux I__2366 (
            .O(N__10860),
            .I(N__10840));
    InMux I__2365 (
            .O(N__10859),
            .I(N__10840));
    Odrv4 I__2364 (
            .O(N__10856),
            .I(buart__rx_bitcount_3));
    LocalMux I__2363 (
            .O(N__10853),
            .I(buart__rx_bitcount_3));
    LocalMux I__2362 (
            .O(N__10850),
            .I(buart__rx_bitcount_3));
    LocalMux I__2361 (
            .O(N__10847),
            .I(buart__rx_bitcount_3));
    LocalMux I__2360 (
            .O(N__10840),
            .I(buart__rx_bitcount_3));
    CascadeMux I__2359 (
            .O(N__10829),
            .I(N__10826));
    InMux I__2358 (
            .O(N__10826),
            .I(N__10822));
    InMux I__2357 (
            .O(N__10825),
            .I(N__10814));
    LocalMux I__2356 (
            .O(N__10822),
            .I(N__10811));
    InMux I__2355 (
            .O(N__10821),
            .I(N__10808));
    InMux I__2354 (
            .O(N__10820),
            .I(N__10799));
    InMux I__2353 (
            .O(N__10819),
            .I(N__10799));
    InMux I__2352 (
            .O(N__10818),
            .I(N__10799));
    InMux I__2351 (
            .O(N__10817),
            .I(N__10799));
    LocalMux I__2350 (
            .O(N__10814),
            .I(buart__rx_bitcount_2));
    Odrv4 I__2349 (
            .O(N__10811),
            .I(buart__rx_bitcount_2));
    LocalMux I__2348 (
            .O(N__10808),
            .I(buart__rx_bitcount_2));
    LocalMux I__2347 (
            .O(N__10799),
            .I(buart__rx_bitcount_2));
    InMux I__2346 (
            .O(N__10790),
            .I(N__10787));
    LocalMux I__2345 (
            .O(N__10787),
            .I(N__10784));
    Span4Mux_v I__2344 (
            .O(N__10784),
            .I(N__10779));
    InMux I__2343 (
            .O(N__10783),
            .I(N__10774));
    InMux I__2342 (
            .O(N__10782),
            .I(N__10774));
    Odrv4 I__2341 (
            .O(N__10779),
            .I(N_87));
    LocalMux I__2340 (
            .O(N__10774),
            .I(N_87));
    InMux I__2339 (
            .O(N__10769),
            .I(N__10766));
    LocalMux I__2338 (
            .O(N__10766),
            .I(\Lab_UT.rx_data_rdy ));
    InMux I__2337 (
            .O(N__10763),
            .I(N__10755));
    InMux I__2336 (
            .O(N__10762),
            .I(N__10755));
    InMux I__2335 (
            .O(N__10761),
            .I(N__10749));
    InMux I__2334 (
            .O(N__10760),
            .I(N__10746));
    LocalMux I__2333 (
            .O(N__10755),
            .I(N__10743));
    InMux I__2332 (
            .O(N__10754),
            .I(N__10740));
    InMux I__2331 (
            .O(N__10753),
            .I(N__10735));
    InMux I__2330 (
            .O(N__10752),
            .I(N__10735));
    LocalMux I__2329 (
            .O(N__10749),
            .I(buart__rx_bitcount_0));
    LocalMux I__2328 (
            .O(N__10746),
            .I(buart__rx_bitcount_0));
    Odrv4 I__2327 (
            .O(N__10743),
            .I(buart__rx_bitcount_0));
    LocalMux I__2326 (
            .O(N__10740),
            .I(buart__rx_bitcount_0));
    LocalMux I__2325 (
            .O(N__10735),
            .I(buart__rx_bitcount_0));
    InMux I__2324 (
            .O(N__10724),
            .I(N__10721));
    LocalMux I__2323 (
            .O(N__10721),
            .I(N__10718));
    Span4Mux_h I__2322 (
            .O(N__10718),
            .I(N__10715));
    Odrv4 I__2321 (
            .O(N__10715),
            .I(\resetGen.un3_reset_count_i_a3Z0Z_4 ));
    InMux I__2320 (
            .O(N__10712),
            .I(N__10709));
    LocalMux I__2319 (
            .O(N__10709),
            .I(N__10706));
    Span4Mux_v I__2318 (
            .O(N__10706),
            .I(N__10703));
    Span4Mux_h I__2317 (
            .O(N__10703),
            .I(N__10700));
    Odrv4 I__2316 (
            .O(N__10700),
            .I(Lab_UT_L3_tx_data_0_6));
    InMux I__2315 (
            .O(N__10697),
            .I(N__10692));
    InMux I__2314 (
            .O(N__10696),
            .I(N__10686));
    InMux I__2313 (
            .O(N__10695),
            .I(N__10686));
    LocalMux I__2312 (
            .O(N__10692),
            .I(N__10683));
    CascadeMux I__2311 (
            .O(N__10691),
            .I(N__10680));
    LocalMux I__2310 (
            .O(N__10686),
            .I(N__10676));
    Span4Mux_v I__2309 (
            .O(N__10683),
            .I(N__10670));
    InMux I__2308 (
            .O(N__10680),
            .I(N__10667));
    InMux I__2307 (
            .O(N__10679),
            .I(N__10661));
    Span4Mux_v I__2306 (
            .O(N__10676),
            .I(N__10658));
    InMux I__2305 (
            .O(N__10675),
            .I(N__10655));
    InMux I__2304 (
            .O(N__10674),
            .I(N__10650));
    InMux I__2303 (
            .O(N__10673),
            .I(N__10650));
    Span4Mux_h I__2302 (
            .O(N__10670),
            .I(N__10645));
    LocalMux I__2301 (
            .O(N__10667),
            .I(N__10645));
    InMux I__2300 (
            .O(N__10666),
            .I(N__10638));
    InMux I__2299 (
            .O(N__10665),
            .I(N__10638));
    InMux I__2298 (
            .O(N__10664),
            .I(N__10638));
    LocalMux I__2297 (
            .O(N__10661),
            .I(Lab_UT_dspStr_cnt_2));
    Odrv4 I__2296 (
            .O(N__10658),
            .I(Lab_UT_dspStr_cnt_2));
    LocalMux I__2295 (
            .O(N__10655),
            .I(Lab_UT_dspStr_cnt_2));
    LocalMux I__2294 (
            .O(N__10650),
            .I(Lab_UT_dspStr_cnt_2));
    Odrv4 I__2293 (
            .O(N__10645),
            .I(Lab_UT_dspStr_cnt_2));
    LocalMux I__2292 (
            .O(N__10638),
            .I(Lab_UT_dspStr_cnt_2));
    CascadeMux I__2291 (
            .O(N__10625),
            .I(N__10621));
    CascadeMux I__2290 (
            .O(N__10624),
            .I(N__10614));
    InMux I__2289 (
            .O(N__10621),
            .I(N__10610));
    CascadeMux I__2288 (
            .O(N__10620),
            .I(N__10607));
    CascadeMux I__2287 (
            .O(N__10619),
            .I(N__10604));
    CascadeMux I__2286 (
            .O(N__10618),
            .I(N__10601));
    InMux I__2285 (
            .O(N__10617),
            .I(N__10596));
    InMux I__2284 (
            .O(N__10614),
            .I(N__10596));
    CascadeMux I__2283 (
            .O(N__10613),
            .I(N__10592));
    LocalMux I__2282 (
            .O(N__10610),
            .I(N__10588));
    InMux I__2281 (
            .O(N__10607),
            .I(N__10583));
    InMux I__2280 (
            .O(N__10604),
            .I(N__10583));
    InMux I__2279 (
            .O(N__10601),
            .I(N__10580));
    LocalMux I__2278 (
            .O(N__10596),
            .I(N__10575));
    InMux I__2277 (
            .O(N__10595),
            .I(N__10568));
    InMux I__2276 (
            .O(N__10592),
            .I(N__10568));
    InMux I__2275 (
            .O(N__10591),
            .I(N__10568));
    Span4Mux_v I__2274 (
            .O(N__10588),
            .I(N__10563));
    LocalMux I__2273 (
            .O(N__10583),
            .I(N__10563));
    LocalMux I__2272 (
            .O(N__10580),
            .I(N__10560));
    InMux I__2271 (
            .O(N__10579),
            .I(N__10557));
    InMux I__2270 (
            .O(N__10578),
            .I(N__10554));
    Span4Mux_v I__2269 (
            .O(N__10575),
            .I(N__10549));
    LocalMux I__2268 (
            .O(N__10568),
            .I(N__10549));
    Span4Mux_h I__2267 (
            .O(N__10563),
            .I(N__10546));
    Span4Mux_h I__2266 (
            .O(N__10560),
            .I(N__10543));
    LocalMux I__2265 (
            .O(N__10557),
            .I(Lab_UT_dspStr_cnt_3));
    LocalMux I__2264 (
            .O(N__10554),
            .I(Lab_UT_dspStr_cnt_3));
    Odrv4 I__2263 (
            .O(N__10549),
            .I(Lab_UT_dspStr_cnt_3));
    Odrv4 I__2262 (
            .O(N__10546),
            .I(Lab_UT_dspStr_cnt_3));
    Odrv4 I__2261 (
            .O(N__10543),
            .I(Lab_UT_dspStr_cnt_3));
    InMux I__2260 (
            .O(N__10532),
            .I(N__10529));
    LocalMux I__2259 (
            .O(N__10529),
            .I(\buart.Z_tx.bitcount_RNO_0Z0Z_2 ));
    InMux I__2258 (
            .O(N__10526),
            .I(\buart.Z_tx.un1_bitcount_cry_1 ));
    CascadeMux I__2257 (
            .O(N__10523),
            .I(N__10520));
    InMux I__2256 (
            .O(N__10520),
            .I(N__10513));
    CascadeMux I__2255 (
            .O(N__10519),
            .I(N__10510));
    InMux I__2254 (
            .O(N__10518),
            .I(N__10500));
    InMux I__2253 (
            .O(N__10517),
            .I(N__10500));
    InMux I__2252 (
            .O(N__10516),
            .I(N__10497));
    LocalMux I__2251 (
            .O(N__10513),
            .I(N__10494));
    InMux I__2250 (
            .O(N__10510),
            .I(N__10489));
    InMux I__2249 (
            .O(N__10509),
            .I(N__10489));
    CascadeMux I__2248 (
            .O(N__10508),
            .I(N__10481));
    CascadeMux I__2247 (
            .O(N__10507),
            .I(N__10478));
    CascadeMux I__2246 (
            .O(N__10506),
            .I(N__10473));
    InMux I__2245 (
            .O(N__10505),
            .I(N__10466));
    LocalMux I__2244 (
            .O(N__10500),
            .I(N__10457));
    LocalMux I__2243 (
            .O(N__10497),
            .I(N__10457));
    Span4Mux_h I__2242 (
            .O(N__10494),
            .I(N__10457));
    LocalMux I__2241 (
            .O(N__10489),
            .I(N__10457));
    InMux I__2240 (
            .O(N__10488),
            .I(N__10450));
    InMux I__2239 (
            .O(N__10487),
            .I(N__10450));
    InMux I__2238 (
            .O(N__10486),
            .I(N__10450));
    InMux I__2237 (
            .O(N__10485),
            .I(N__10445));
    InMux I__2236 (
            .O(N__10484),
            .I(N__10445));
    InMux I__2235 (
            .O(N__10481),
            .I(N__10438));
    InMux I__2234 (
            .O(N__10478),
            .I(N__10438));
    InMux I__2233 (
            .O(N__10477),
            .I(N__10438));
    InMux I__2232 (
            .O(N__10476),
            .I(N__10431));
    InMux I__2231 (
            .O(N__10473),
            .I(N__10431));
    InMux I__2230 (
            .O(N__10472),
            .I(N__10431));
    InMux I__2229 (
            .O(N__10471),
            .I(N__10424));
    InMux I__2228 (
            .O(N__10470),
            .I(N__10424));
    InMux I__2227 (
            .O(N__10469),
            .I(N__10424));
    LocalMux I__2226 (
            .O(N__10466),
            .I(N__10421));
    Span4Mux_h I__2225 (
            .O(N__10457),
            .I(N__10418));
    LocalMux I__2224 (
            .O(N__10450),
            .I(uu2_un3_r_clk_en_0));
    LocalMux I__2223 (
            .O(N__10445),
            .I(uu2_un3_r_clk_en_0));
    LocalMux I__2222 (
            .O(N__10438),
            .I(uu2_un3_r_clk_en_0));
    LocalMux I__2221 (
            .O(N__10431),
            .I(uu2_un3_r_clk_en_0));
    LocalMux I__2220 (
            .O(N__10424),
            .I(uu2_un3_r_clk_en_0));
    Odrv12 I__2219 (
            .O(N__10421),
            .I(uu2_un3_r_clk_en_0));
    Odrv4 I__2218 (
            .O(N__10418),
            .I(uu2_un3_r_clk_en_0));
    InMux I__2217 (
            .O(N__10403),
            .I(\buart.Z_tx.un1_bitcount_cry_2 ));
    InMux I__2216 (
            .O(N__10400),
            .I(N__10397));
    LocalMux I__2215 (
            .O(N__10397),
            .I(\buart.Z_tx.bitcount_RNIM5O32Z0Z_2 ));
    CascadeMux I__2214 (
            .O(N__10394),
            .I(N__10390));
    InMux I__2213 (
            .O(N__10393),
            .I(N__10384));
    InMux I__2212 (
            .O(N__10390),
            .I(N__10384));
    InMux I__2211 (
            .O(N__10389),
            .I(N__10381));
    LocalMux I__2210 (
            .O(N__10384),
            .I(N__10376));
    LocalMux I__2209 (
            .O(N__10381),
            .I(N__10376));
    Odrv4 I__2208 (
            .O(N__10376),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__2207 (
            .O(N__10373),
            .I(N__10368));
    InMux I__2206 (
            .O(N__10372),
            .I(N__10362));
    InMux I__2205 (
            .O(N__10371),
            .I(N__10362));
    InMux I__2204 (
            .O(N__10368),
            .I(N__10357));
    InMux I__2203 (
            .O(N__10367),
            .I(N__10357));
    LocalMux I__2202 (
            .O(N__10362),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__2201 (
            .O(N__10357),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    CascadeMux I__2200 (
            .O(N__10352),
            .I(N__10349));
    InMux I__2199 (
            .O(N__10349),
            .I(N__10344));
    InMux I__2198 (
            .O(N__10348),
            .I(N__10339));
    InMux I__2197 (
            .O(N__10347),
            .I(N__10339));
    LocalMux I__2196 (
            .O(N__10344),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    LocalMux I__2195 (
            .O(N__10339),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    CascadeMux I__2194 (
            .O(N__10334),
            .I(buart__tx_uart_busy_0_cascade_));
    InMux I__2193 (
            .O(N__10331),
            .I(N__10328));
    LocalMux I__2192 (
            .O(N__10328),
            .I(\buart.Z_tx.bitcount_RNIL4O32Z0Z_1 ));
    InMux I__2191 (
            .O(N__10325),
            .I(N__10310));
    InMux I__2190 (
            .O(N__10324),
            .I(N__10310));
    InMux I__2189 (
            .O(N__10323),
            .I(N__10310));
    InMux I__2188 (
            .O(N__10322),
            .I(N__10303));
    InMux I__2187 (
            .O(N__10321),
            .I(N__10303));
    InMux I__2186 (
            .O(N__10320),
            .I(N__10303));
    InMux I__2185 (
            .O(N__10319),
            .I(N__10296));
    InMux I__2184 (
            .O(N__10318),
            .I(N__10296));
    InMux I__2183 (
            .O(N__10317),
            .I(N__10296));
    LocalMux I__2182 (
            .O(N__10310),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__2181 (
            .O(N__10303),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__2180 (
            .O(N__10296),
            .I(\buart.Z_tx.ser_clk ));
    CascadeMux I__2179 (
            .O(N__10289),
            .I(N__10281));
    InMux I__2178 (
            .O(N__10288),
            .I(N__10265));
    InMux I__2177 (
            .O(N__10287),
            .I(N__10265));
    InMux I__2176 (
            .O(N__10286),
            .I(N__10265));
    InMux I__2175 (
            .O(N__10285),
            .I(N__10265));
    CascadeMux I__2174 (
            .O(N__10284),
            .I(N__10262));
    InMux I__2173 (
            .O(N__10281),
            .I(N__10259));
    InMux I__2172 (
            .O(N__10280),
            .I(N__10254));
    InMux I__2171 (
            .O(N__10279),
            .I(N__10254));
    InMux I__2170 (
            .O(N__10278),
            .I(N__10245));
    InMux I__2169 (
            .O(N__10277),
            .I(N__10245));
    InMux I__2168 (
            .O(N__10276),
            .I(N__10245));
    InMux I__2167 (
            .O(N__10275),
            .I(N__10245));
    CascadeMux I__2166 (
            .O(N__10274),
            .I(N__10241));
    LocalMux I__2165 (
            .O(N__10265),
            .I(N__10233));
    InMux I__2164 (
            .O(N__10262),
            .I(N__10230));
    LocalMux I__2163 (
            .O(N__10259),
            .I(N__10223));
    LocalMux I__2162 (
            .O(N__10254),
            .I(N__10223));
    LocalMux I__2161 (
            .O(N__10245),
            .I(N__10223));
    InMux I__2160 (
            .O(N__10244),
            .I(N__10216));
    InMux I__2159 (
            .O(N__10241),
            .I(N__10216));
    InMux I__2158 (
            .O(N__10240),
            .I(N__10216));
    InMux I__2157 (
            .O(N__10239),
            .I(N__10207));
    InMux I__2156 (
            .O(N__10238),
            .I(N__10207));
    InMux I__2155 (
            .O(N__10237),
            .I(N__10207));
    InMux I__2154 (
            .O(N__10236),
            .I(N__10207));
    Span4Mux_h I__2153 (
            .O(N__10233),
            .I(N__10204));
    LocalMux I__2152 (
            .O(N__10230),
            .I(buart__tx_uart_busy_0));
    Odrv4 I__2151 (
            .O(N__10223),
            .I(buart__tx_uart_busy_0));
    LocalMux I__2150 (
            .O(N__10216),
            .I(buart__tx_uart_busy_0));
    LocalMux I__2149 (
            .O(N__10207),
            .I(buart__tx_uart_busy_0));
    Odrv4 I__2148 (
            .O(N__10204),
            .I(buart__tx_uart_busy_0));
    CascadeMux I__2147 (
            .O(N__10193),
            .I(N__10189));
    InMux I__2146 (
            .O(N__10192),
            .I(N__10186));
    InMux I__2145 (
            .O(N__10189),
            .I(N__10183));
    LocalMux I__2144 (
            .O(N__10186),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    LocalMux I__2143 (
            .O(N__10183),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    InMux I__2142 (
            .O(N__10178),
            .I(N__10175));
    LocalMux I__2141 (
            .O(N__10175),
            .I(\buart.Z_tx.un1_bitcount_axb_3 ));
    CascadeMux I__2140 (
            .O(N__10172),
            .I(N__10169));
    InMux I__2139 (
            .O(N__10169),
            .I(N__10165));
    InMux I__2138 (
            .O(N__10168),
            .I(N__10162));
    LocalMux I__2137 (
            .O(N__10165),
            .I(N__10159));
    LocalMux I__2136 (
            .O(N__10162),
            .I(\Lab_UT.dspStr.cnt11_0_i ));
    Odrv4 I__2135 (
            .O(N__10159),
            .I(\Lab_UT.dspStr.cnt11_0_i ));
    InMux I__2134 (
            .O(N__10154),
            .I(N__10151));
    LocalMux I__2133 (
            .O(N__10151),
            .I(N__10148));
    Span4Mux_v I__2132 (
            .O(N__10148),
            .I(N__10145));
    Span4Mux_h I__2131 (
            .O(N__10145),
            .I(N__10140));
    InMux I__2130 (
            .O(N__10144),
            .I(N__10137));
    InMux I__2129 (
            .O(N__10143),
            .I(N__10134));
    Odrv4 I__2128 (
            .O(N__10140),
            .I(\Lab_UT.dspStr.cntZ0Z_0 ));
    LocalMux I__2127 (
            .O(N__10137),
            .I(\Lab_UT.dspStr.cntZ0Z_0 ));
    LocalMux I__2126 (
            .O(N__10134),
            .I(\Lab_UT.dspStr.cntZ0Z_0 ));
    InMux I__2125 (
            .O(N__10127),
            .I(\Lab_UT.didpuu0.didpsones.un1_q_cry_0 ));
    InMux I__2124 (
            .O(N__10124),
            .I(N__10121));
    LocalMux I__2123 (
            .O(N__10121),
            .I(\Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_2 ));
    InMux I__2122 (
            .O(N__10118),
            .I(\Lab_UT.didpuu0.didpsones.un1_q_cry_1 ));
    InMux I__2121 (
            .O(N__10115),
            .I(\Lab_UT.didpuu0.didpsones.un1_q_cry_2 ));
    CascadeMux I__2120 (
            .O(N__10112),
            .I(\Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_3_cascade_ ));
    InMux I__2119 (
            .O(N__10109),
            .I(N__10106));
    LocalMux I__2118 (
            .O(N__10106),
            .I(\Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_0 ));
    InMux I__2117 (
            .O(N__10103),
            .I(N__10100));
    LocalMux I__2116 (
            .O(N__10100),
            .I(\Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_1 ));
    CascadeMux I__2115 (
            .O(N__10097),
            .I(N__10092));
    CascadeMux I__2114 (
            .O(N__10096),
            .I(N__10089));
    InMux I__2113 (
            .O(N__10095),
            .I(N__10082));
    InMux I__2112 (
            .O(N__10092),
            .I(N__10082));
    InMux I__2111 (
            .O(N__10089),
            .I(N__10082));
    LocalMux I__2110 (
            .O(N__10082),
            .I(\Lab_UT.didpuu0.didpsones.q13_0 ));
    InMux I__2109 (
            .O(N__10079),
            .I(N__10069));
    InMux I__2108 (
            .O(N__10078),
            .I(N__10069));
    InMux I__2107 (
            .O(N__10077),
            .I(N__10069));
    InMux I__2106 (
            .O(N__10076),
            .I(N__10066));
    LocalMux I__2105 (
            .O(N__10069),
            .I(N__10060));
    LocalMux I__2104 (
            .O(N__10066),
            .I(N__10060));
    InMux I__2103 (
            .O(N__10065),
            .I(N__10056));
    Span4Mux_h I__2102 (
            .O(N__10060),
            .I(N__10053));
    InMux I__2101 (
            .O(N__10059),
            .I(N__10050));
    LocalMux I__2100 (
            .O(N__10056),
            .I(N__10047));
    Span4Mux_v I__2099 (
            .O(N__10053),
            .I(N__10044));
    LocalMux I__2098 (
            .O(N__10050),
            .I(N__10039));
    Span4Mux_h I__2097 (
            .O(N__10047),
            .I(N__10039));
    Odrv4 I__2096 (
            .O(N__10044),
            .I(rst));
    Odrv4 I__2095 (
            .O(N__10039),
            .I(rst));
    InMux I__2094 (
            .O(N__10034),
            .I(N__10031));
    LocalMux I__2093 (
            .O(N__10031),
            .I(\buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0 ));
    InMux I__2092 (
            .O(N__10028),
            .I(N__10025));
    LocalMux I__2091 (
            .O(N__10025),
            .I(\buart.Z_tx.bitcount_RNO_0Z0Z_1 ));
    InMux I__2090 (
            .O(N__10022),
            .I(\buart.Z_tx.un1_bitcount_cry_0 ));
    CascadeMux I__2089 (
            .O(N__10019),
            .I(N__10015));
    CascadeMux I__2088 (
            .O(N__10018),
            .I(N__10011));
    InMux I__2087 (
            .O(N__10015),
            .I(N__10008));
    InMux I__2086 (
            .O(N__10014),
            .I(N__10002));
    InMux I__2085 (
            .O(N__10011),
            .I(N__9999));
    LocalMux I__2084 (
            .O(N__10008),
            .I(N__9996));
    InMux I__2083 (
            .O(N__10007),
            .I(N__9989));
    InMux I__2082 (
            .O(N__10006),
            .I(N__9989));
    InMux I__2081 (
            .O(N__10005),
            .I(N__9989));
    LocalMux I__2080 (
            .O(N__10002),
            .I(\uu2.w_addr_displaying_fastZ0Z_4 ));
    LocalMux I__2079 (
            .O(N__9999),
            .I(\uu2.w_addr_displaying_fastZ0Z_4 ));
    Odrv4 I__2078 (
            .O(N__9996),
            .I(\uu2.w_addr_displaying_fastZ0Z_4 ));
    LocalMux I__2077 (
            .O(N__9989),
            .I(\uu2.w_addr_displaying_fastZ0Z_4 ));
    InMux I__2076 (
            .O(N__9980),
            .I(N__9977));
    LocalMux I__2075 (
            .O(N__9977),
            .I(N__9974));
    Odrv4 I__2074 (
            .O(N__9974),
            .I(\uu2.mem0.Z_decfrac105_7_3_2 ));
    CascadeMux I__2073 (
            .O(N__9971),
            .I(\uu2.w_addr_displaying_4_8_cascade_ ));
    CascadeMux I__2072 (
            .O(N__9968),
            .I(N__9961));
    InMux I__2071 (
            .O(N__9967),
            .I(N__9958));
    CascadeMux I__2070 (
            .O(N__9966),
            .I(N__9954));
    InMux I__2069 (
            .O(N__9965),
            .I(N__9951));
    InMux I__2068 (
            .O(N__9964),
            .I(N__9946));
    InMux I__2067 (
            .O(N__9961),
            .I(N__9946));
    LocalMux I__2066 (
            .O(N__9958),
            .I(N__9940));
    InMux I__2065 (
            .O(N__9957),
            .I(N__9937));
    InMux I__2064 (
            .O(N__9954),
            .I(N__9934));
    LocalMux I__2063 (
            .O(N__9951),
            .I(N__9929));
    LocalMux I__2062 (
            .O(N__9946),
            .I(N__9929));
    InMux I__2061 (
            .O(N__9945),
            .I(N__9922));
    InMux I__2060 (
            .O(N__9944),
            .I(N__9922));
    InMux I__2059 (
            .O(N__9943),
            .I(N__9922));
    Span4Mux_h I__2058 (
            .O(N__9940),
            .I(N__9917));
    LocalMux I__2057 (
            .O(N__9937),
            .I(N__9917));
    LocalMux I__2056 (
            .O(N__9934),
            .I(N__9914));
    Span4Mux_v I__2055 (
            .O(N__9929),
            .I(N__9911));
    LocalMux I__2054 (
            .O(N__9922),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2053 (
            .O(N__9917),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2052 (
            .O(N__9914),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2051 (
            .O(N__9911),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    InMux I__2050 (
            .O(N__9902),
            .I(N__9896));
    InMux I__2049 (
            .O(N__9901),
            .I(N__9893));
    InMux I__2048 (
            .O(N__9900),
            .I(N__9888));
    InMux I__2047 (
            .O(N__9899),
            .I(N__9888));
    LocalMux I__2046 (
            .O(N__9896),
            .I(N__9885));
    LocalMux I__2045 (
            .O(N__9893),
            .I(N__9880));
    LocalMux I__2044 (
            .O(N__9888),
            .I(N__9880));
    Odrv12 I__2043 (
            .O(N__9885),
            .I(\uu2.un15_w_data_displaying ));
    Odrv4 I__2042 (
            .O(N__9880),
            .I(\uu2.un15_w_data_displaying ));
    CascadeMux I__2041 (
            .O(N__9875),
            .I(\uu2.un15_w_data_displaying_cascade_ ));
    CascadeMux I__2040 (
            .O(N__9872),
            .I(N__9866));
    CascadeMux I__2039 (
            .O(N__9871),
            .I(N__9862));
    InMux I__2038 (
            .O(N__9870),
            .I(N__9858));
    InMux I__2037 (
            .O(N__9869),
            .I(N__9855));
    InMux I__2036 (
            .O(N__9866),
            .I(N__9852));
    InMux I__2035 (
            .O(N__9865),
            .I(N__9849));
    InMux I__2034 (
            .O(N__9862),
            .I(N__9844));
    InMux I__2033 (
            .O(N__9861),
            .I(N__9844));
    LocalMux I__2032 (
            .O(N__9858),
            .I(N__9839));
    LocalMux I__2031 (
            .O(N__9855),
            .I(N__9834));
    LocalMux I__2030 (
            .O(N__9852),
            .I(N__9834));
    LocalMux I__2029 (
            .O(N__9849),
            .I(N__9829));
    LocalMux I__2028 (
            .O(N__9844),
            .I(N__9829));
    InMux I__2027 (
            .O(N__9843),
            .I(N__9826));
    InMux I__2026 (
            .O(N__9842),
            .I(N__9823));
    Span4Mux_v I__2025 (
            .O(N__9839),
            .I(N__9820));
    Span4Mux_v I__2024 (
            .O(N__9834),
            .I(N__9817));
    Span4Mux_v I__2023 (
            .O(N__9829),
            .I(N__9814));
    LocalMux I__2022 (
            .O(N__9826),
            .I(N__9811));
    LocalMux I__2021 (
            .O(N__9823),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2020 (
            .O(N__9820),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2019 (
            .O(N__9817),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2018 (
            .O(N__9814),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2017 (
            .O(N__9811),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    InMux I__2016 (
            .O(N__9800),
            .I(N__9797));
    LocalMux I__2015 (
            .O(N__9797),
            .I(N__9792));
    InMux I__2014 (
            .O(N__9796),
            .I(N__9789));
    InMux I__2013 (
            .O(N__9795),
            .I(N__9784));
    Span4Mux_h I__2012 (
            .O(N__9792),
            .I(N__9781));
    LocalMux I__2011 (
            .O(N__9789),
            .I(N__9778));
    InMux I__2010 (
            .O(N__9788),
            .I(N__9773));
    InMux I__2009 (
            .O(N__9787),
            .I(N__9773));
    LocalMux I__2008 (
            .O(N__9784),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    Odrv4 I__2007 (
            .O(N__9781),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    Odrv4 I__2006 (
            .O(N__9778),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__2005 (
            .O(N__9773),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    CascadeMux I__2004 (
            .O(N__9764),
            .I(N__9757));
    CascadeMux I__2003 (
            .O(N__9763),
            .I(N__9754));
    CascadeMux I__2002 (
            .O(N__9762),
            .I(N__9751));
    CascadeMux I__2001 (
            .O(N__9761),
            .I(N__9746));
    CascadeMux I__2000 (
            .O(N__9760),
            .I(N__9743));
    InMux I__1999 (
            .O(N__9757),
            .I(N__9738));
    InMux I__1998 (
            .O(N__9754),
            .I(N__9738));
    InMux I__1997 (
            .O(N__9751),
            .I(N__9731));
    InMux I__1996 (
            .O(N__9750),
            .I(N__9731));
    InMux I__1995 (
            .O(N__9749),
            .I(N__9731));
    InMux I__1994 (
            .O(N__9746),
            .I(N__9726));
    InMux I__1993 (
            .O(N__9743),
            .I(N__9726));
    LocalMux I__1992 (
            .O(N__9738),
            .I(N__9723));
    LocalMux I__1991 (
            .O(N__9731),
            .I(N__9718));
    LocalMux I__1990 (
            .O(N__9726),
            .I(N__9718));
    Span4Mux_v I__1989 (
            .O(N__9723),
            .I(N__9715));
    Span4Mux_v I__1988 (
            .O(N__9718),
            .I(N__9712));
    Odrv4 I__1987 (
            .O(N__9715),
            .I(\uu2.un448_ci_5 ));
    Odrv4 I__1986 (
            .O(N__9712),
            .I(\uu2.un448_ci_5 ));
    InMux I__1985 (
            .O(N__9707),
            .I(N__9700));
    InMux I__1984 (
            .O(N__9706),
            .I(N__9696));
    InMux I__1983 (
            .O(N__9705),
            .I(N__9692));
    InMux I__1982 (
            .O(N__9704),
            .I(N__9689));
    CascadeMux I__1981 (
            .O(N__9703),
            .I(N__9685));
    LocalMux I__1980 (
            .O(N__9700),
            .I(N__9682));
    InMux I__1979 (
            .O(N__9699),
            .I(N__9679));
    LocalMux I__1978 (
            .O(N__9696),
            .I(N__9676));
    InMux I__1977 (
            .O(N__9695),
            .I(N__9673));
    LocalMux I__1976 (
            .O(N__9692),
            .I(N__9664));
    LocalMux I__1975 (
            .O(N__9689),
            .I(N__9664));
    InMux I__1974 (
            .O(N__9688),
            .I(N__9659));
    InMux I__1973 (
            .O(N__9685),
            .I(N__9659));
    Span4Mux_v I__1972 (
            .O(N__9682),
            .I(N__9654));
    LocalMux I__1971 (
            .O(N__9679),
            .I(N__9654));
    Span4Mux_v I__1970 (
            .O(N__9676),
            .I(N__9649));
    LocalMux I__1969 (
            .O(N__9673),
            .I(N__9649));
    InMux I__1968 (
            .O(N__9672),
            .I(N__9640));
    InMux I__1967 (
            .O(N__9671),
            .I(N__9640));
    InMux I__1966 (
            .O(N__9670),
            .I(N__9640));
    InMux I__1965 (
            .O(N__9669),
            .I(N__9640));
    Span4Mux_v I__1964 (
            .O(N__9664),
            .I(N__9637));
    LocalMux I__1963 (
            .O(N__9659),
            .I(N__9634));
    Span4Mux_h I__1962 (
            .O(N__9654),
            .I(N__9631));
    Span4Mux_v I__1961 (
            .O(N__9649),
            .I(N__9628));
    LocalMux I__1960 (
            .O(N__9640),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__1959 (
            .O(N__9637),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__1958 (
            .O(N__9634),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__1957 (
            .O(N__9631),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__1956 (
            .O(N__9628),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    InMux I__1955 (
            .O(N__9617),
            .I(N__9608));
    InMux I__1954 (
            .O(N__9616),
            .I(N__9608));
    InMux I__1953 (
            .O(N__9615),
            .I(N__9608));
    LocalMux I__1952 (
            .O(N__9608),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    InMux I__1951 (
            .O(N__9605),
            .I(N__9599));
    InMux I__1950 (
            .O(N__9604),
            .I(N__9590));
    InMux I__1949 (
            .O(N__9603),
            .I(N__9590));
    InMux I__1948 (
            .O(N__9602),
            .I(N__9590));
    LocalMux I__1947 (
            .O(N__9599),
            .I(N__9586));
    InMux I__1946 (
            .O(N__9598),
            .I(N__9583));
    InMux I__1945 (
            .O(N__9597),
            .I(N__9578));
    LocalMux I__1944 (
            .O(N__9590),
            .I(N__9575));
    InMux I__1943 (
            .O(N__9589),
            .I(N__9572));
    Span4Mux_v I__1942 (
            .O(N__9586),
            .I(N__9567));
    LocalMux I__1941 (
            .O(N__9583),
            .I(N__9567));
    InMux I__1940 (
            .O(N__9582),
            .I(N__9564));
    InMux I__1939 (
            .O(N__9581),
            .I(N__9561));
    LocalMux I__1938 (
            .O(N__9578),
            .I(N__9556));
    Span4Mux_h I__1937 (
            .O(N__9575),
            .I(N__9556));
    LocalMux I__1936 (
            .O(N__9572),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    Odrv4 I__1935 (
            .O(N__9567),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    LocalMux I__1934 (
            .O(N__9564),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    LocalMux I__1933 (
            .O(N__9561),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    Odrv4 I__1932 (
            .O(N__9556),
            .I(\uu2.w_addr_displaying_6_repZ0Z1 ));
    InMux I__1931 (
            .O(N__9545),
            .I(N__9541));
    CascadeMux I__1930 (
            .O(N__9544),
            .I(N__9535));
    LocalMux I__1929 (
            .O(N__9541),
            .I(N__9531));
    InMux I__1928 (
            .O(N__9540),
            .I(N__9528));
    CascadeMux I__1927 (
            .O(N__9539),
            .I(N__9524));
    InMux I__1926 (
            .O(N__9538),
            .I(N__9519));
    InMux I__1925 (
            .O(N__9535),
            .I(N__9516));
    InMux I__1924 (
            .O(N__9534),
            .I(N__9513));
    Span4Mux_h I__1923 (
            .O(N__9531),
            .I(N__9510));
    LocalMux I__1922 (
            .O(N__9528),
            .I(N__9507));
    InMux I__1921 (
            .O(N__9527),
            .I(N__9504));
    InMux I__1920 (
            .O(N__9524),
            .I(N__9497));
    InMux I__1919 (
            .O(N__9523),
            .I(N__9497));
    InMux I__1918 (
            .O(N__9522),
            .I(N__9497));
    LocalMux I__1917 (
            .O(N__9519),
            .I(N__9494));
    LocalMux I__1916 (
            .O(N__9516),
            .I(N__9489));
    LocalMux I__1915 (
            .O(N__9513),
            .I(N__9489));
    Odrv4 I__1914 (
            .O(N__9510),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    Odrv4 I__1913 (
            .O(N__9507),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    LocalMux I__1912 (
            .O(N__9504),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    LocalMux I__1911 (
            .O(N__9497),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    Odrv4 I__1910 (
            .O(N__9494),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    Odrv4 I__1909 (
            .O(N__9489),
            .I(\uu2.w_addr_displaying_5_repZ0Z1 ));
    InMux I__1908 (
            .O(N__9476),
            .I(N__9473));
    LocalMux I__1907 (
            .O(N__9473),
            .I(\uu2.mem0.bitmap_pmux_1_1_i_a5_1_0 ));
    CascadeMux I__1906 (
            .O(N__9470),
            .I(\uu2.mem0.g1_1_0_cascade_ ));
    InMux I__1905 (
            .O(N__9467),
            .I(N__9464));
    LocalMux I__1904 (
            .O(N__9464),
            .I(N__9459));
    InMux I__1903 (
            .O(N__9463),
            .I(N__9456));
    InMux I__1902 (
            .O(N__9462),
            .I(N__9453));
    Span4Mux_h I__1901 (
            .O(N__9459),
            .I(N__9448));
    LocalMux I__1900 (
            .O(N__9456),
            .I(N__9448));
    LocalMux I__1899 (
            .O(N__9453),
            .I(N__9445));
    Odrv4 I__1898 (
            .O(N__9448),
            .I(\uu2.Z_decfrac106_5 ));
    Odrv4 I__1897 (
            .O(N__9445),
            .I(\uu2.Z_decfrac106_5 ));
    InMux I__1896 (
            .O(N__9440),
            .I(N__9437));
    LocalMux I__1895 (
            .O(N__9437),
            .I(N__9434));
    Span12Mux_s7_h I__1894 (
            .O(N__9434),
            .I(N__9431));
    Odrv12 I__1893 (
            .O(N__9431),
            .I(\uu2.mem0.g0_2_0 ));
    InMux I__1892 (
            .O(N__9428),
            .I(N__9425));
    LocalMux I__1891 (
            .O(N__9425),
            .I(\uu2.mem0.bitmap_pmux_1_1_i_a5_2_3_1_0 ));
    InMux I__1890 (
            .O(N__9422),
            .I(N__9416));
    CascadeMux I__1889 (
            .O(N__9421),
            .I(N__9413));
    InMux I__1888 (
            .O(N__9420),
            .I(N__9406));
    InMux I__1887 (
            .O(N__9419),
            .I(N__9403));
    LocalMux I__1886 (
            .O(N__9416),
            .I(N__9400));
    InMux I__1885 (
            .O(N__9413),
            .I(N__9397));
    InMux I__1884 (
            .O(N__9412),
            .I(N__9392));
    InMux I__1883 (
            .O(N__9411),
            .I(N__9392));
    InMux I__1882 (
            .O(N__9410),
            .I(N__9389));
    InMux I__1881 (
            .O(N__9409),
            .I(N__9386));
    LocalMux I__1880 (
            .O(N__9406),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__1879 (
            .O(N__9403),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    Odrv4 I__1878 (
            .O(N__9400),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__1877 (
            .O(N__9397),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__1876 (
            .O(N__9392),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__1875 (
            .O(N__9389),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__1874 (
            .O(N__9386),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    InMux I__1873 (
            .O(N__9371),
            .I(N__9362));
    InMux I__1872 (
            .O(N__9370),
            .I(N__9362));
    InMux I__1871 (
            .O(N__9369),
            .I(N__9362));
    LocalMux I__1870 (
            .O(N__9362),
            .I(N__9358));
    InMux I__1869 (
            .O(N__9361),
            .I(N__9355));
    Span4Mux_h I__1868 (
            .O(N__9358),
            .I(N__9352));
    LocalMux I__1867 (
            .O(N__9355),
            .I(N__9349));
    Odrv4 I__1866 (
            .O(N__9352),
            .I(\uu2.Z_decfrac105_7_2 ));
    Odrv4 I__1865 (
            .O(N__9349),
            .I(\uu2.Z_decfrac105_7_2 ));
    CascadeMux I__1864 (
            .O(N__9344),
            .I(N__9339));
    InMux I__1863 (
            .O(N__9343),
            .I(N__9331));
    InMux I__1862 (
            .O(N__9342),
            .I(N__9331));
    InMux I__1861 (
            .O(N__9339),
            .I(N__9331));
    InMux I__1860 (
            .O(N__9338),
            .I(N__9328));
    LocalMux I__1859 (
            .O(N__9331),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    LocalMux I__1858 (
            .O(N__9328),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    CascadeMux I__1857 (
            .O(N__9323),
            .I(L3_tx_data_0_cascade_));
    InMux I__1856 (
            .O(N__9320),
            .I(N__9317));
    LocalMux I__1855 (
            .O(N__9317),
            .I(N__9314));
    Span4Mux_h I__1854 (
            .O(N__9314),
            .I(N__9308));
    InMux I__1853 (
            .O(N__9313),
            .I(N__9301));
    InMux I__1852 (
            .O(N__9312),
            .I(N__9301));
    InMux I__1851 (
            .O(N__9311),
            .I(N__9301));
    Odrv4 I__1850 (
            .O(N__9308),
            .I(\uu2.un1_w_user_crZ0Z_1 ));
    LocalMux I__1849 (
            .O(N__9301),
            .I(\uu2.un1_w_user_crZ0Z_1 ));
    CascadeMux I__1848 (
            .O(N__9296),
            .I(\uu2.w_addr_displaying_RNIQKOV8Z0Z_8_cascade_ ));
    InMux I__1847 (
            .O(N__9293),
            .I(N__9281));
    InMux I__1846 (
            .O(N__9292),
            .I(N__9281));
    InMux I__1845 (
            .O(N__9291),
            .I(N__9281));
    InMux I__1844 (
            .O(N__9290),
            .I(N__9281));
    LocalMux I__1843 (
            .O(N__9281),
            .I(N__9276));
    InMux I__1842 (
            .O(N__9280),
            .I(N__9273));
    InMux I__1841 (
            .O(N__9279),
            .I(N__9270));
    Span4Mux_h I__1840 (
            .O(N__9276),
            .I(N__9267));
    LocalMux I__1839 (
            .O(N__9273),
            .I(L3_tx_data_rdy));
    LocalMux I__1838 (
            .O(N__9270),
            .I(L3_tx_data_rdy));
    Odrv4 I__1837 (
            .O(N__9267),
            .I(L3_tx_data_rdy));
    CascadeMux I__1836 (
            .O(N__9260),
            .I(\uu2.un21_w_addr_displaying_i_cascade_ ));
    CascadeMux I__1835 (
            .O(N__9257),
            .I(N__9254));
    InMux I__1834 (
            .O(N__9254),
            .I(N__9251));
    LocalMux I__1833 (
            .O(N__9251),
            .I(N__9248));
    Span4Mux_h I__1832 (
            .O(N__9248),
            .I(N__9245));
    Odrv4 I__1831 (
            .O(N__9245),
            .I(\uu2.mem0.g0_i_a11_1_0 ));
    CascadeMux I__1830 (
            .O(N__9242),
            .I(N__9239));
    InMux I__1829 (
            .O(N__9239),
            .I(N__9232));
    InMux I__1828 (
            .O(N__9238),
            .I(N__9229));
    InMux I__1827 (
            .O(N__9237),
            .I(N__9225));
    InMux I__1826 (
            .O(N__9236),
            .I(N__9220));
    InMux I__1825 (
            .O(N__9235),
            .I(N__9220));
    LocalMux I__1824 (
            .O(N__9232),
            .I(N__9217));
    LocalMux I__1823 (
            .O(N__9229),
            .I(N__9214));
    CascadeMux I__1822 (
            .O(N__9228),
            .I(N__9211));
    LocalMux I__1821 (
            .O(N__9225),
            .I(N__9206));
    LocalMux I__1820 (
            .O(N__9220),
            .I(N__9199));
    Span4Mux_h I__1819 (
            .O(N__9217),
            .I(N__9199));
    Span4Mux_h I__1818 (
            .O(N__9214),
            .I(N__9196));
    InMux I__1817 (
            .O(N__9211),
            .I(N__9193));
    InMux I__1816 (
            .O(N__9210),
            .I(N__9188));
    InMux I__1815 (
            .O(N__9209),
            .I(N__9188));
    Span4Mux_v I__1814 (
            .O(N__9206),
            .I(N__9185));
    InMux I__1813 (
            .O(N__9205),
            .I(N__9180));
    InMux I__1812 (
            .O(N__9204),
            .I(N__9180));
    Odrv4 I__1811 (
            .O(N__9199),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    Odrv4 I__1810 (
            .O(N__9196),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    LocalMux I__1809 (
            .O(N__9193),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    LocalMux I__1808 (
            .O(N__9188),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    Odrv4 I__1807 (
            .O(N__9185),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    LocalMux I__1806 (
            .O(N__9180),
            .I(\uu2.w_addr_displaying_4_repZ0Z1 ));
    CascadeMux I__1805 (
            .O(N__9167),
            .I(\uu2.mem0.g3_0_cascade_ ));
    InMux I__1804 (
            .O(N__9164),
            .I(N__9157));
    InMux I__1803 (
            .O(N__9163),
            .I(N__9157));
    InMux I__1802 (
            .O(N__9162),
            .I(N__9152));
    LocalMux I__1801 (
            .O(N__9157),
            .I(N__9149));
    InMux I__1800 (
            .O(N__9156),
            .I(N__9145));
    InMux I__1799 (
            .O(N__9155),
            .I(N__9142));
    LocalMux I__1798 (
            .O(N__9152),
            .I(N__9139));
    Span4Mux_v I__1797 (
            .O(N__9149),
            .I(N__9129));
    InMux I__1796 (
            .O(N__9148),
            .I(N__9126));
    LocalMux I__1795 (
            .O(N__9145),
            .I(N__9123));
    LocalMux I__1794 (
            .O(N__9142),
            .I(N__9120));
    Span4Mux_h I__1793 (
            .O(N__9139),
            .I(N__9117));
    InMux I__1792 (
            .O(N__9138),
            .I(N__9110));
    InMux I__1791 (
            .O(N__9137),
            .I(N__9110));
    InMux I__1790 (
            .O(N__9136),
            .I(N__9110));
    InMux I__1789 (
            .O(N__9135),
            .I(N__9103));
    InMux I__1788 (
            .O(N__9134),
            .I(N__9103));
    InMux I__1787 (
            .O(N__9133),
            .I(N__9103));
    InMux I__1786 (
            .O(N__9132),
            .I(N__9100));
    Odrv4 I__1785 (
            .O(N__9129),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__1784 (
            .O(N__9126),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__1783 (
            .O(N__9123),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__1782 (
            .O(N__9120),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__1781 (
            .O(N__9117),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__1780 (
            .O(N__9110),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__1779 (
            .O(N__9103),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__1778 (
            .O(N__9100),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    InMux I__1777 (
            .O(N__9083),
            .I(N__9080));
    LocalMux I__1776 (
            .O(N__9080),
            .I(N__9077));
    Odrv4 I__1775 (
            .O(N__9077),
            .I(\uu2.mem0.un1_segment4_0_i_i_0_0 ));
    InMux I__1774 (
            .O(N__9074),
            .I(N__9071));
    LocalMux I__1773 (
            .O(N__9071),
            .I(N__9068));
    Odrv12 I__1772 (
            .O(N__9068),
            .I(\uu2.mem0.g0_i_a11_3_1 ));
    CascadeMux I__1771 (
            .O(N__9065),
            .I(\uu2.mem0.g0_i_a11_7_1_cascade_ ));
    InMux I__1770 (
            .O(N__9062),
            .I(N__9059));
    LocalMux I__1769 (
            .O(N__9059),
            .I(N__9056));
    Odrv4 I__1768 (
            .O(N__9056),
            .I(\uu2.mem0.g0_i_5_1 ));
    InMux I__1767 (
            .O(N__9053),
            .I(N__9047));
    InMux I__1766 (
            .O(N__9052),
            .I(N__9040));
    InMux I__1765 (
            .O(N__9051),
            .I(N__9040));
    InMux I__1764 (
            .O(N__9050),
            .I(N__9040));
    LocalMux I__1763 (
            .O(N__9047),
            .I(Lab_UT_dspStr_cnt_1_rep1));
    LocalMux I__1762 (
            .O(N__9040),
            .I(Lab_UT_dspStr_cnt_1_rep1));
    InMux I__1761 (
            .O(N__9035),
            .I(N__9032));
    LocalMux I__1760 (
            .O(N__9032),
            .I(N__9029));
    Span4Mux_h I__1759 (
            .O(N__9029),
            .I(N__9026));
    Odrv4 I__1758 (
            .O(N__9026),
            .I(Lab_UT_dspStr_un36_dOut));
    CascadeMux I__1757 (
            .O(N__9023),
            .I(Lab_UT_dspStr_un36_dOut_cascade_));
    CascadeMux I__1756 (
            .O(N__9020),
            .I(\uu2.un27_N_6_mux_cascade_ ));
    InMux I__1755 (
            .O(N__9017),
            .I(N__9014));
    LocalMux I__1754 (
            .O(N__9014),
            .I(N__9011));
    Odrv4 I__1753 (
            .O(N__9011),
            .I(\uu2.un27_w_addr_user_iZ0Z_1 ));
    CascadeMux I__1752 (
            .O(N__9008),
            .I(N__9003));
    CascadeMux I__1751 (
            .O(N__9007),
            .I(N__9000));
    InMux I__1750 (
            .O(N__9006),
            .I(N__8996));
    InMux I__1749 (
            .O(N__9003),
            .I(N__8989));
    InMux I__1748 (
            .O(N__9000),
            .I(N__8989));
    InMux I__1747 (
            .O(N__8999),
            .I(N__8989));
    LocalMux I__1746 (
            .O(N__8996),
            .I(Lab_UT_dspStr_cnt_3_rep1));
    LocalMux I__1745 (
            .O(N__8989),
            .I(Lab_UT_dspStr_cnt_3_rep1));
    InMux I__1744 (
            .O(N__8984),
            .I(N__8975));
    InMux I__1743 (
            .O(N__8983),
            .I(N__8975));
    InMux I__1742 (
            .O(N__8982),
            .I(N__8968));
    InMux I__1741 (
            .O(N__8981),
            .I(N__8968));
    InMux I__1740 (
            .O(N__8980),
            .I(N__8968));
    LocalMux I__1739 (
            .O(N__8975),
            .I(Lab_UT_dspStr_cnt_2_rep1));
    LocalMux I__1738 (
            .O(N__8968),
            .I(Lab_UT_dspStr_cnt_2_rep1));
    InMux I__1737 (
            .O(N__8963),
            .I(N__8960));
    LocalMux I__1736 (
            .O(N__8960),
            .I(N__8956));
    CascadeMux I__1735 (
            .O(N__8959),
            .I(N__8953));
    Span4Mux_h I__1734 (
            .O(N__8956),
            .I(N__8950));
    InMux I__1733 (
            .O(N__8953),
            .I(N__8947));
    Odrv4 I__1732 (
            .O(N__8950),
            .I(L3_tx_data_0));
    LocalMux I__1731 (
            .O(N__8947),
            .I(L3_tx_data_0));
    InMux I__1730 (
            .O(N__8942),
            .I(N__8939));
    LocalMux I__1729 (
            .O(N__8939),
            .I(\uu2.w_m5_i_a3Z0Z_2 ));
    InMux I__1728 (
            .O(N__8936),
            .I(N__8933));
    LocalMux I__1727 (
            .O(N__8933),
            .I(\Lab_UT.dictrluu0.dek.det_NZ0Z_4 ));
    CascadeMux I__1726 (
            .O(N__8930),
            .I(\uu2.un1_w_user_lf_0_0Z0Z_0_cascade_ ));
    InMux I__1725 (
            .O(N__8927),
            .I(N__8924));
    LocalMux I__1724 (
            .O(N__8924),
            .I(\uu2.un1_w_user_lf_2 ));
    InMux I__1723 (
            .O(N__8921),
            .I(N__8918));
    LocalMux I__1722 (
            .O(N__8918),
            .I(N__8914));
    InMux I__1721 (
            .O(N__8917),
            .I(N__8911));
    Span4Mux_v I__1720 (
            .O(N__8914),
            .I(N__8908));
    LocalMux I__1719 (
            .O(N__8911),
            .I(\uu2.un2_w_addr_user ));
    Odrv4 I__1718 (
            .O(N__8908),
            .I(\uu2.un2_w_addr_user ));
    CascadeMux I__1717 (
            .O(N__8903),
            .I(\uu2.un1_w_user_lf_2_cascade_ ));
    InMux I__1716 (
            .O(N__8900),
            .I(N__8897));
    LocalMux I__1715 (
            .O(N__8897),
            .I(\uu2.un27_N_6_mux_0 ));
    IoInMux I__1714 (
            .O(N__8894),
            .I(N__8889));
    InMux I__1713 (
            .O(N__8893),
            .I(N__8886));
    CascadeMux I__1712 (
            .O(N__8892),
            .I(N__8883));
    LocalMux I__1711 (
            .O(N__8889),
            .I(N__8880));
    LocalMux I__1710 (
            .O(N__8886),
            .I(N__8877));
    InMux I__1709 (
            .O(N__8883),
            .I(N__8874));
    Span4Mux_s2_v I__1708 (
            .O(N__8880),
            .I(N__8871));
    Span4Mux_h I__1707 (
            .O(N__8877),
            .I(N__8866));
    LocalMux I__1706 (
            .O(N__8874),
            .I(N__8866));
    Span4Mux_h I__1705 (
            .O(N__8871),
            .I(N__8863));
    Odrv4 I__1704 (
            .O(N__8866),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1703 (
            .O(N__8863),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1702 (
            .O(N__8858),
            .I(\uu2.w_addr_user_RNILDNK6Z0Z_4_cascade_ ));
    InMux I__1701 (
            .O(N__8855),
            .I(N__8848));
    InMux I__1700 (
            .O(N__8854),
            .I(N__8848));
    InMux I__1699 (
            .O(N__8853),
            .I(N__8839));
    LocalMux I__1698 (
            .O(N__8848),
            .I(N__8836));
    InMux I__1697 (
            .O(N__8847),
            .I(N__8829));
    InMux I__1696 (
            .O(N__8846),
            .I(N__8829));
    InMux I__1695 (
            .O(N__8845),
            .I(N__8829));
    InMux I__1694 (
            .O(N__8844),
            .I(N__8822));
    InMux I__1693 (
            .O(N__8843),
            .I(N__8822));
    InMux I__1692 (
            .O(N__8842),
            .I(N__8822));
    LocalMux I__1691 (
            .O(N__8839),
            .I(N__8819));
    Odrv4 I__1690 (
            .O(N__8836),
            .I(\uu2.un27_w_addr_user_i ));
    LocalMux I__1689 (
            .O(N__8829),
            .I(\uu2.un27_w_addr_user_i ));
    LocalMux I__1688 (
            .O(N__8822),
            .I(\uu2.un27_w_addr_user_i ));
    Odrv4 I__1687 (
            .O(N__8819),
            .I(\uu2.un27_w_addr_user_i ));
    CascadeMux I__1686 (
            .O(N__8810),
            .I(\uu2.un1_w_user_lf_5_a0Z0Z_5_cascade_ ));
    InMux I__1685 (
            .O(N__8807),
            .I(N__8804));
    LocalMux I__1684 (
            .O(N__8804),
            .I(N__8800));
    InMux I__1683 (
            .O(N__8803),
            .I(N__8797));
    Odrv4 I__1682 (
            .O(N__8800),
            .I(\uu2.un1_w_user_lf_5_aZ0Z0 ));
    LocalMux I__1681 (
            .O(N__8797),
            .I(\uu2.un1_w_user_lf_5_aZ0Z0 ));
    CascadeMux I__1680 (
            .O(N__8792),
            .I(\uu2.w_addr_user_2Z0Z_1_cascade_ ));
    CascadeMux I__1679 (
            .O(N__8789),
            .I(\uu2.w_addr_userZ2Z_1_cascade_ ));
    SRMux I__1678 (
            .O(N__8786),
            .I(N__8782));
    SRMux I__1677 (
            .O(N__8785),
            .I(N__8778));
    LocalMux I__1676 (
            .O(N__8782),
            .I(N__8774));
    SRMux I__1675 (
            .O(N__8781),
            .I(N__8771));
    LocalMux I__1674 (
            .O(N__8778),
            .I(N__8768));
    SRMux I__1673 (
            .O(N__8777),
            .I(N__8765));
    Span4Mux_h I__1672 (
            .O(N__8774),
            .I(N__8762));
    LocalMux I__1671 (
            .O(N__8771),
            .I(N__8755));
    Span4Mux_s3_v I__1670 (
            .O(N__8768),
            .I(N__8755));
    LocalMux I__1669 (
            .O(N__8765),
            .I(N__8755));
    Odrv4 I__1668 (
            .O(N__8762),
            .I(\uu2.w_addr_user_RNIT1MGDZ0Z_4 ));
    Odrv4 I__1667 (
            .O(N__8755),
            .I(\uu2.w_addr_user_RNIT1MGDZ0Z_4 ));
    InMux I__1666 (
            .O(N__8750),
            .I(N__8747));
    LocalMux I__1665 (
            .O(N__8747),
            .I(\uu2.w_addr_user_1_0 ));
    CascadeMux I__1664 (
            .O(N__8744),
            .I(\Lab_UT.dictrluu0.dek.det_NZ0Z_5_cascade_ ));
    InMux I__1663 (
            .O(N__8741),
            .I(N__8738));
    LocalMux I__1662 (
            .O(N__8738),
            .I(N__8735));
    Span4Mux_v I__1661 (
            .O(N__8735),
            .I(N__8732));
    Odrv4 I__1660 (
            .O(N__8732),
            .I(\uu2.mem0.N_1476_0_0_0 ));
    InMux I__1659 (
            .O(N__8729),
            .I(N__8726));
    LocalMux I__1658 (
            .O(N__8726),
            .I(\Lab_UT.dspStr.cnt11_1 ));
    InMux I__1657 (
            .O(N__8723),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__1656 (
            .O(N__8720),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__1655 (
            .O(N__8717),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__1654 (
            .O(N__8714),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__1653 (
            .O(N__8711),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    CascadeMux I__1652 (
            .O(N__8708),
            .I(N__8705));
    InMux I__1651 (
            .O(N__8705),
            .I(N__8699));
    InMux I__1650 (
            .O(N__8704),
            .I(N__8699));
    LocalMux I__1649 (
            .O(N__8699),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__1648 (
            .O(N__8696),
            .I(N__8693));
    InMux I__1647 (
            .O(N__8693),
            .I(N__8687));
    InMux I__1646 (
            .O(N__8692),
            .I(N__8687));
    LocalMux I__1645 (
            .O(N__8687),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__1644 (
            .O(N__8684),
            .I(N__8680));
    InMux I__1643 (
            .O(N__8683),
            .I(N__8677));
    InMux I__1642 (
            .O(N__8680),
            .I(N__8674));
    LocalMux I__1641 (
            .O(N__8677),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    LocalMux I__1640 (
            .O(N__8674),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    InMux I__1639 (
            .O(N__8669),
            .I(N__8663));
    InMux I__1638 (
            .O(N__8668),
            .I(N__8663));
    LocalMux I__1637 (
            .O(N__8663),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    CascadeMux I__1636 (
            .O(N__8660),
            .I(N__8656));
    InMux I__1635 (
            .O(N__8659),
            .I(N__8652));
    InMux I__1634 (
            .O(N__8656),
            .I(N__8649));
    InMux I__1633 (
            .O(N__8655),
            .I(N__8646));
    LocalMux I__1632 (
            .O(N__8652),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1631 (
            .O(N__8649),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1630 (
            .O(N__8646),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    InMux I__1629 (
            .O(N__8639),
            .I(N__8631));
    InMux I__1628 (
            .O(N__8638),
            .I(N__8631));
    InMux I__1627 (
            .O(N__8637),
            .I(N__8628));
    InMux I__1626 (
            .O(N__8636),
            .I(N__8625));
    LocalMux I__1625 (
            .O(N__8631),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1624 (
            .O(N__8628),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1623 (
            .O(N__8625),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__1622 (
            .O(N__8618),
            .I(N__8614));
    CascadeMux I__1621 (
            .O(N__8617),
            .I(N__8611));
    InMux I__1620 (
            .O(N__8614),
            .I(N__8606));
    InMux I__1619 (
            .O(N__8611),
            .I(N__8606));
    LocalMux I__1618 (
            .O(N__8606),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    InMux I__1617 (
            .O(N__8603),
            .I(N__8600));
    LocalMux I__1616 (
            .O(N__8600),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    CascadeMux I__1615 (
            .O(N__8597),
            .I(\Lab_UT.didpuu0.didpsones.q13_0_cascade_ ));
    InMux I__1614 (
            .O(N__8594),
            .I(N__8591));
    LocalMux I__1613 (
            .O(N__8591),
            .I(\uu2.g0_3Z0Z_0 ));
    CEMux I__1612 (
            .O(N__8588),
            .I(N__8585));
    LocalMux I__1611 (
            .O(N__8585),
            .I(N__8580));
    CEMux I__1610 (
            .O(N__8584),
            .I(N__8577));
    CEMux I__1609 (
            .O(N__8583),
            .I(N__8574));
    Span4Mux_v I__1608 (
            .O(N__8580),
            .I(N__8571));
    LocalMux I__1607 (
            .O(N__8577),
            .I(N__8568));
    LocalMux I__1606 (
            .O(N__8574),
            .I(N__8565));
    Span4Mux_h I__1605 (
            .O(N__8571),
            .I(N__8562));
    Span4Mux_h I__1604 (
            .O(N__8568),
            .I(N__8559));
    Span4Mux_h I__1603 (
            .O(N__8565),
            .I(N__8556));
    Odrv4 I__1602 (
            .O(N__8562),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__1601 (
            .O(N__8559),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__1600 (
            .O(N__8556),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    InMux I__1599 (
            .O(N__8549),
            .I(N__8543));
    InMux I__1598 (
            .O(N__8548),
            .I(N__8538));
    InMux I__1597 (
            .O(N__8547),
            .I(N__8538));
    InMux I__1596 (
            .O(N__8546),
            .I(N__8535));
    LocalMux I__1595 (
            .O(N__8543),
            .I(N__8529));
    LocalMux I__1594 (
            .O(N__8538),
            .I(N__8529));
    LocalMux I__1593 (
            .O(N__8535),
            .I(N__8526));
    CascadeMux I__1592 (
            .O(N__8534),
            .I(N__8522));
    Span4Mux_h I__1591 (
            .O(N__8529),
            .I(N__8517));
    Span4Mux_h I__1590 (
            .O(N__8526),
            .I(N__8514));
    InMux I__1589 (
            .O(N__8525),
            .I(N__8511));
    InMux I__1588 (
            .O(N__8522),
            .I(N__8506));
    InMux I__1587 (
            .O(N__8521),
            .I(N__8506));
    InMux I__1586 (
            .O(N__8520),
            .I(N__8503));
    Odrv4 I__1585 (
            .O(N__8517),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    Odrv4 I__1584 (
            .O(N__8514),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__1583 (
            .O(N__8511),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__1582 (
            .O(N__8506),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__1581 (
            .O(N__8503),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    InMux I__1580 (
            .O(N__8492),
            .I(N__8489));
    LocalMux I__1579 (
            .O(N__8489),
            .I(N__8486));
    Span4Mux_h I__1578 (
            .O(N__8486),
            .I(N__8483));
    Odrv4 I__1577 (
            .O(N__8483),
            .I(\uu2.mem0.N_10_0 ));
    CascadeMux I__1576 (
            .O(N__8480),
            .I(\uu2.w_addr_displaying_4_rep1_3_cascade_ ));
    CascadeMux I__1575 (
            .O(N__8477),
            .I(N__8474));
    InMux I__1574 (
            .O(N__8474),
            .I(N__8468));
    InMux I__1573 (
            .O(N__8473),
            .I(N__8468));
    LocalMux I__1572 (
            .O(N__8468),
            .I(N__8463));
    InMux I__1571 (
            .O(N__8467),
            .I(N__8456));
    InMux I__1570 (
            .O(N__8466),
            .I(N__8456));
    Span4Mux_h I__1569 (
            .O(N__8463),
            .I(N__8453));
    InMux I__1568 (
            .O(N__8462),
            .I(N__8448));
    InMux I__1567 (
            .O(N__8461),
            .I(N__8448));
    LocalMux I__1566 (
            .O(N__8456),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    Odrv4 I__1565 (
            .O(N__8453),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__1564 (
            .O(N__8448),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    CascadeMux I__1563 (
            .O(N__8441),
            .I(N__8438));
    InMux I__1562 (
            .O(N__8438),
            .I(N__8432));
    InMux I__1561 (
            .O(N__8437),
            .I(N__8432));
    LocalMux I__1560 (
            .O(N__8432),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    InMux I__1559 (
            .O(N__8429),
            .I(N__8426));
    LocalMux I__1558 (
            .O(N__8426),
            .I(\uu2.mem0.un1_segment4_0_i_i_1 ));
    InMux I__1557 (
            .O(N__8423),
            .I(N__8420));
    LocalMux I__1556 (
            .O(N__8420),
            .I(\uu2.mem0.un1_segment4_0_i_i_a5_0_0 ));
    InMux I__1555 (
            .O(N__8417),
            .I(N__8413));
    InMux I__1554 (
            .O(N__8416),
            .I(N__8410));
    LocalMux I__1553 (
            .O(N__8413),
            .I(N__8403));
    LocalMux I__1552 (
            .O(N__8410),
            .I(N__8400));
    CascadeMux I__1551 (
            .O(N__8409),
            .I(N__8393));
    InMux I__1550 (
            .O(N__8408),
            .I(N__8390));
    InMux I__1549 (
            .O(N__8407),
            .I(N__8387));
    InMux I__1548 (
            .O(N__8406),
            .I(N__8384));
    Span4Mux_h I__1547 (
            .O(N__8403),
            .I(N__8381));
    Span4Mux_h I__1546 (
            .O(N__8400),
            .I(N__8378));
    InMux I__1545 (
            .O(N__8399),
            .I(N__8375));
    InMux I__1544 (
            .O(N__8398),
            .I(N__8366));
    InMux I__1543 (
            .O(N__8397),
            .I(N__8366));
    InMux I__1542 (
            .O(N__8396),
            .I(N__8366));
    InMux I__1541 (
            .O(N__8393),
            .I(N__8366));
    LocalMux I__1540 (
            .O(N__8390),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__1539 (
            .O(N__8387),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__1538 (
            .O(N__8384),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    Odrv4 I__1537 (
            .O(N__8381),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    Odrv4 I__1536 (
            .O(N__8378),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__1535 (
            .O(N__8375),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__1534 (
            .O(N__8366),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    CascadeMux I__1533 (
            .O(N__8351),
            .I(\uu2.g1_0_1_cascade_ ));
    CascadeMux I__1532 (
            .O(N__8348),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_50_cascade_ ));
    InMux I__1531 (
            .O(N__8345),
            .I(N__8342));
    LocalMux I__1530 (
            .O(N__8342),
            .I(\uu2.g1_0_1 ));
    InMux I__1529 (
            .O(N__8339),
            .I(N__8336));
    LocalMux I__1528 (
            .O(N__8336),
            .I(\uu2.mem0.g0_0 ));
    InMux I__1527 (
            .O(N__8333),
            .I(N__8329));
    InMux I__1526 (
            .O(N__8332),
            .I(N__8325));
    LocalMux I__1525 (
            .O(N__8329),
            .I(N__8321));
    InMux I__1524 (
            .O(N__8328),
            .I(N__8318));
    LocalMux I__1523 (
            .O(N__8325),
            .I(N__8315));
    InMux I__1522 (
            .O(N__8324),
            .I(N__8305));
    Span4Mux_v I__1521 (
            .O(N__8321),
            .I(N__8302));
    LocalMux I__1520 (
            .O(N__8318),
            .I(N__8297));
    Span4Mux_h I__1519 (
            .O(N__8315),
            .I(N__8297));
    InMux I__1518 (
            .O(N__8314),
            .I(N__8292));
    InMux I__1517 (
            .O(N__8313),
            .I(N__8292));
    InMux I__1516 (
            .O(N__8312),
            .I(N__8287));
    InMux I__1515 (
            .O(N__8311),
            .I(N__8287));
    InMux I__1514 (
            .O(N__8310),
            .I(N__8280));
    InMux I__1513 (
            .O(N__8309),
            .I(N__8280));
    InMux I__1512 (
            .O(N__8308),
            .I(N__8280));
    LocalMux I__1511 (
            .O(N__8305),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    Odrv4 I__1510 (
            .O(N__8302),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    Odrv4 I__1509 (
            .O(N__8297),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    LocalMux I__1508 (
            .O(N__8292),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    LocalMux I__1507 (
            .O(N__8287),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    LocalMux I__1506 (
            .O(N__8280),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    CascadeMux I__1505 (
            .O(N__8267),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_ ));
    CascadeMux I__1504 (
            .O(N__8264),
            .I(N__8261));
    InMux I__1503 (
            .O(N__8261),
            .I(N__8258));
    LocalMux I__1502 (
            .O(N__8258),
            .I(N__8255));
    Odrv4 I__1501 (
            .O(N__8255),
            .I(\uu2.mem0.g1 ));
    InMux I__1500 (
            .O(N__8252),
            .I(N__8243));
    InMux I__1499 (
            .O(N__8251),
            .I(N__8243));
    InMux I__1498 (
            .O(N__8250),
            .I(N__8243));
    LocalMux I__1497 (
            .O(N__8243),
            .I(\uu2.N_10 ));
    InMux I__1496 (
            .O(N__8240),
            .I(N__8237));
    LocalMux I__1495 (
            .O(N__8237),
            .I(\uu2.mem0.g1_1_1 ));
    CascadeMux I__1494 (
            .O(N__8234),
            .I(\uu2.mem0.w_data_ns_1_1_0_3_cascade_ ));
    InMux I__1493 (
            .O(N__8231),
            .I(N__8224));
    InMux I__1492 (
            .O(N__8230),
            .I(N__8224));
    InMux I__1491 (
            .O(N__8229),
            .I(N__8221));
    LocalMux I__1490 (
            .O(N__8224),
            .I(\uu2.Z_decfrac106 ));
    LocalMux I__1489 (
            .O(N__8221),
            .I(\uu2.Z_decfrac106 ));
    InMux I__1488 (
            .O(N__8216),
            .I(N__8213));
    LocalMux I__1487 (
            .O(N__8213),
            .I(\uu2.mem0.w_data_ns_1_0_0_1_3 ));
    CascadeMux I__1486 (
            .O(N__8210),
            .I(\uu2.g0_1_0_0_1_cascade_ ));
    InMux I__1485 (
            .O(N__8207),
            .I(N__8201));
    InMux I__1484 (
            .O(N__8206),
            .I(N__8201));
    LocalMux I__1483 (
            .O(N__8201),
            .I(\uu2.g0_1_0_0 ));
    CascadeMux I__1482 (
            .O(N__8198),
            .I(N__8195));
    InMux I__1481 (
            .O(N__8195),
            .I(N__8192));
    LocalMux I__1480 (
            .O(N__8192),
            .I(\uu2.g0_1_a5_0_0 ));
    InMux I__1479 (
            .O(N__8189),
            .I(N__8186));
    LocalMux I__1478 (
            .O(N__8186),
            .I(N__8183));
    Odrv4 I__1477 (
            .O(N__8183),
            .I(\uu2.g0_1_a5_1_0 ));
    InMux I__1476 (
            .O(N__8180),
            .I(N__8174));
    InMux I__1475 (
            .O(N__8179),
            .I(N__8174));
    LocalMux I__1474 (
            .O(N__8174),
            .I(\uu2.g1_1 ));
    InMux I__1473 (
            .O(N__8171),
            .I(N__8168));
    LocalMux I__1472 (
            .O(N__8168),
            .I(N__8162));
    InMux I__1471 (
            .O(N__8167),
            .I(N__8159));
    InMux I__1470 (
            .O(N__8166),
            .I(N__8154));
    InMux I__1469 (
            .O(N__8165),
            .I(N__8154));
    Span4Mux_h I__1468 (
            .O(N__8162),
            .I(N__8151));
    LocalMux I__1467 (
            .O(N__8159),
            .I(N__8148));
    LocalMux I__1466 (
            .O(N__8154),
            .I(\uu2.w_addr_userZ0Z_8 ));
    Odrv4 I__1465 (
            .O(N__8151),
            .I(\uu2.w_addr_userZ0Z_8 ));
    Odrv4 I__1464 (
            .O(N__8148),
            .I(\uu2.w_addr_userZ0Z_8 ));
    InMux I__1463 (
            .O(N__8141),
            .I(N__8128));
    InMux I__1462 (
            .O(N__8140),
            .I(N__8128));
    InMux I__1461 (
            .O(N__8139),
            .I(N__8128));
    InMux I__1460 (
            .O(N__8138),
            .I(N__8128));
    InMux I__1459 (
            .O(N__8137),
            .I(N__8125));
    LocalMux I__1458 (
            .O(N__8128),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__1457 (
            .O(N__8125),
            .I(\uu2.w_addr_userZ0Z_7 ));
    InMux I__1456 (
            .O(N__8120),
            .I(N__8116));
    CascadeMux I__1455 (
            .O(N__8119),
            .I(N__8112));
    LocalMux I__1454 (
            .O(N__8116),
            .I(N__8107));
    InMux I__1453 (
            .O(N__8115),
            .I(N__8104));
    InMux I__1452 (
            .O(N__8112),
            .I(N__8097));
    InMux I__1451 (
            .O(N__8111),
            .I(N__8097));
    InMux I__1450 (
            .O(N__8110),
            .I(N__8097));
    Span4Mux_h I__1449 (
            .O(N__8107),
            .I(N__8092));
    LocalMux I__1448 (
            .O(N__8104),
            .I(N__8092));
    LocalMux I__1447 (
            .O(N__8097),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv4 I__1446 (
            .O(N__8092),
            .I(\uu2.w_addr_userZ0Z_2 ));
    InMux I__1445 (
            .O(N__8087),
            .I(N__8082));
    CascadeMux I__1444 (
            .O(N__8086),
            .I(N__8078));
    CascadeMux I__1443 (
            .O(N__8085),
            .I(N__8075));
    LocalMux I__1442 (
            .O(N__8082),
            .I(N__8071));
    InMux I__1441 (
            .O(N__8081),
            .I(N__8068));
    InMux I__1440 (
            .O(N__8078),
            .I(N__8061));
    InMux I__1439 (
            .O(N__8075),
            .I(N__8061));
    InMux I__1438 (
            .O(N__8074),
            .I(N__8061));
    Span4Mux_v I__1437 (
            .O(N__8071),
            .I(N__8058));
    LocalMux I__1436 (
            .O(N__8068),
            .I(N__8055));
    LocalMux I__1435 (
            .O(N__8061),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__1434 (
            .O(N__8058),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__1433 (
            .O(N__8055),
            .I(\uu2.w_addr_userZ0Z_6 ));
    CascadeMux I__1432 (
            .O(N__8048),
            .I(\uu2.un2_w_addr_user_4_cascade_ ));
    InMux I__1431 (
            .O(N__8045),
            .I(N__8042));
    LocalMux I__1430 (
            .O(N__8042),
            .I(N__8039));
    Odrv4 I__1429 (
            .O(N__8039),
            .I(\uu2.un2_w_addr_user_5 ));
    CascadeMux I__1428 (
            .O(N__8036),
            .I(\uu2.un448_ci_5_cascade_ ));
    CascadeMux I__1427 (
            .O(N__8033),
            .I(N__8028));
    CascadeMux I__1426 (
            .O(N__8032),
            .I(N__8025));
    CascadeMux I__1425 (
            .O(N__8031),
            .I(N__8022));
    InMux I__1424 (
            .O(N__8028),
            .I(N__8018));
    InMux I__1423 (
            .O(N__8025),
            .I(N__8015));
    InMux I__1422 (
            .O(N__8022),
            .I(N__8010));
    InMux I__1421 (
            .O(N__8021),
            .I(N__8010));
    LocalMux I__1420 (
            .O(N__8018),
            .I(N__8007));
    LocalMux I__1419 (
            .O(N__8015),
            .I(N__8004));
    LocalMux I__1418 (
            .O(N__8010),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__1417 (
            .O(N__8007),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv12 I__1416 (
            .O(N__8004),
            .I(\uu2.w_addr_userZ0Z_5 ));
    InMux I__1415 (
            .O(N__7997),
            .I(N__7991));
    InMux I__1414 (
            .O(N__7996),
            .I(N__7991));
    LocalMux I__1413 (
            .O(N__7991),
            .I(N__7988));
    Span4Mux_v I__1412 (
            .O(N__7988),
            .I(N__7982));
    InMux I__1411 (
            .O(N__7987),
            .I(N__7975));
    InMux I__1410 (
            .O(N__7986),
            .I(N__7975));
    InMux I__1409 (
            .O(N__7985),
            .I(N__7975));
    Odrv4 I__1408 (
            .O(N__7982),
            .I(\uu2.un415_ci ));
    LocalMux I__1407 (
            .O(N__7975),
            .I(\uu2.un415_ci ));
    InMux I__1406 (
            .O(N__7970),
            .I(N__7963));
    InMux I__1405 (
            .O(N__7969),
            .I(N__7954));
    InMux I__1404 (
            .O(N__7968),
            .I(N__7954));
    InMux I__1403 (
            .O(N__7967),
            .I(N__7954));
    InMux I__1402 (
            .O(N__7966),
            .I(N__7954));
    LocalMux I__1401 (
            .O(N__7963),
            .I(\uu2.w_addr_userZ0Z_4 ));
    LocalMux I__1400 (
            .O(N__7954),
            .I(\uu2.w_addr_userZ0Z_4 ));
    CascadeMux I__1399 (
            .O(N__7949),
            .I(N__7946));
    InMux I__1398 (
            .O(N__7946),
            .I(N__7943));
    LocalMux I__1397 (
            .O(N__7943),
            .I(N__7940));
    Odrv12 I__1396 (
            .O(N__7940),
            .I(\uu2.mem0.w_addr_4 ));
    CascadeMux I__1395 (
            .O(N__7937),
            .I(\uu2.mem0.g0_8_0_cascade_ ));
    InMux I__1394 (
            .O(N__7934),
            .I(N__7931));
    LocalMux I__1393 (
            .O(N__7931),
            .I(N__7924));
    InMux I__1392 (
            .O(N__7930),
            .I(N__7914));
    InMux I__1391 (
            .O(N__7929),
            .I(N__7914));
    InMux I__1390 (
            .O(N__7928),
            .I(N__7914));
    InMux I__1389 (
            .O(N__7927),
            .I(N__7914));
    Span4Mux_h I__1388 (
            .O(N__7924),
            .I(N__7911));
    InMux I__1387 (
            .O(N__7923),
            .I(N__7908));
    LocalMux I__1386 (
            .O(N__7914),
            .I(\uu2.w_addr_userZ1Z_1 ));
    Odrv4 I__1385 (
            .O(N__7911),
            .I(\uu2.w_addr_userZ1Z_1 ));
    LocalMux I__1384 (
            .O(N__7908),
            .I(\uu2.w_addr_userZ1Z_1 ));
    CascadeMux I__1383 (
            .O(N__7901),
            .I(\uu2.o_adder_vbuf_w_addr_user_7_cascade_ ));
    CascadeMux I__1382 (
            .O(N__7898),
            .I(N__7895));
    InMux I__1381 (
            .O(N__7895),
            .I(N__7892));
    LocalMux I__1380 (
            .O(N__7892),
            .I(N__7889));
    Span4Mux_v I__1379 (
            .O(N__7889),
            .I(N__7886));
    Odrv4 I__1378 (
            .O(N__7886),
            .I(\uu2.mem0.w_addr_7 ));
    CascadeMux I__1377 (
            .O(N__7883),
            .I(\uu2.vbuf_w_addr_user.un459_ci_0_cascade_ ));
    CascadeMux I__1376 (
            .O(N__7880),
            .I(\uu2.o_adder_vbuf_w_addr_user_8_cascade_ ));
    InMux I__1375 (
            .O(N__7877),
            .I(N__7870));
    InMux I__1374 (
            .O(N__7876),
            .I(N__7870));
    InMux I__1373 (
            .O(N__7875),
            .I(N__7867));
    LocalMux I__1372 (
            .O(N__7870),
            .I(N__7864));
    LocalMux I__1371 (
            .O(N__7867),
            .I(\uu2.un437_ci_3 ));
    Odrv4 I__1370 (
            .O(N__7864),
            .I(\uu2.un437_ci_3 ));
    InMux I__1369 (
            .O(N__7859),
            .I(N__7855));
    InMux I__1368 (
            .O(N__7858),
            .I(N__7852));
    LocalMux I__1367 (
            .O(N__7855),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    LocalMux I__1366 (
            .O(N__7852),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    InMux I__1365 (
            .O(N__7847),
            .I(N__7844));
    LocalMux I__1364 (
            .O(N__7844),
            .I(vbuf_tx_data_0));
    InMux I__1363 (
            .O(N__7841),
            .I(N__7838));
    LocalMux I__1362 (
            .O(N__7838),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__1361 (
            .O(N__7835),
            .I(N__7832));
    LocalMux I__1360 (
            .O(N__7832),
            .I(vbuf_tx_data_1));
    CascadeMux I__1359 (
            .O(N__7829),
            .I(N__7826));
    InMux I__1358 (
            .O(N__7826),
            .I(N__7823));
    LocalMux I__1357 (
            .O(N__7823),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    CascadeMux I__1356 (
            .O(N__7820),
            .I(N__7817));
    InMux I__1355 (
            .O(N__7817),
            .I(N__7814));
    LocalMux I__1354 (
            .O(N__7814),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    CascadeMux I__1353 (
            .O(N__7811),
            .I(\uu2.o_adder_vbuf_w_addr_user_3_cascade_ ));
    InMux I__1352 (
            .O(N__7808),
            .I(N__7805));
    LocalMux I__1351 (
            .O(N__7805),
            .I(N__7800));
    CascadeMux I__1350 (
            .O(N__7804),
            .I(N__7796));
    CascadeMux I__1349 (
            .O(N__7803),
            .I(N__7793));
    Span4Mux_v I__1348 (
            .O(N__7800),
            .I(N__7789));
    InMux I__1347 (
            .O(N__7799),
            .I(N__7780));
    InMux I__1346 (
            .O(N__7796),
            .I(N__7780));
    InMux I__1345 (
            .O(N__7793),
            .I(N__7780));
    InMux I__1344 (
            .O(N__7792),
            .I(N__7780));
    Odrv4 I__1343 (
            .O(N__7789),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__1342 (
            .O(N__7780),
            .I(\uu2.w_addr_userZ0Z_3 ));
    CascadeMux I__1341 (
            .O(N__7775),
            .I(led_c_0_4_cascade_));
    InMux I__1340 (
            .O(N__7772),
            .I(N__7769));
    LocalMux I__1339 (
            .O(N__7769),
            .I(\uu2.mem0.g1_0_0_0 ));
    CascadeMux I__1338 (
            .O(N__7766),
            .I(N__7763));
    InMux I__1337 (
            .O(N__7763),
            .I(N__7760));
    LocalMux I__1336 (
            .O(N__7760),
            .I(\uu2.mem0.g0_i_5_1_0 ));
    InMux I__1335 (
            .O(N__7757),
            .I(N__7754));
    LocalMux I__1334 (
            .O(N__7754),
            .I(\uu2.mem0.g2_0 ));
    CascadeMux I__1333 (
            .O(N__7751),
            .I(\uu2.w_addr_displaying_4_rep1_8_cascade_ ));
    CascadeMux I__1332 (
            .O(N__7748),
            .I(\uu2.N_42_0_0_cascade_ ));
    CascadeMux I__1331 (
            .O(N__7745),
            .I(N__7742));
    InMux I__1330 (
            .O(N__7742),
            .I(N__7736));
    InMux I__1329 (
            .O(N__7741),
            .I(N__7736));
    LocalMux I__1328 (
            .O(N__7736),
            .I(N__7733));
    Odrv4 I__1327 (
            .O(N__7733),
            .I(\uu2.N_1482_0_0 ));
    CascadeMux I__1326 (
            .O(N__7730),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_34_cascade_ ));
    CascadeMux I__1325 (
            .O(N__7727),
            .I(\uu2.mem0.un1_segment3_m6_0_0_0_0_cascade_ ));
    InMux I__1324 (
            .O(N__7724),
            .I(N__7721));
    LocalMux I__1323 (
            .O(N__7721),
            .I(N__7718));
    Span4Mux_h I__1322 (
            .O(N__7718),
            .I(N__7715));
    Odrv4 I__1321 (
            .O(N__7715),
            .I(\uu2.mem0.w_data_3 ));
    InMux I__1320 (
            .O(N__7712),
            .I(N__7709));
    LocalMux I__1319 (
            .O(N__7709),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_35 ));
    InMux I__1318 (
            .O(N__7706),
            .I(N__7703));
    LocalMux I__1317 (
            .O(N__7703),
            .I(N__7700));
    Odrv12 I__1316 (
            .O(N__7700),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_21 ));
    InMux I__1315 (
            .O(N__7697),
            .I(N__7694));
    LocalMux I__1314 (
            .O(N__7694),
            .I(N__7691));
    Odrv4 I__1313 (
            .O(N__7691),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_22 ));
    InMux I__1312 (
            .O(N__7688),
            .I(N__7685));
    LocalMux I__1311 (
            .O(N__7685),
            .I(N__7682));
    Sp12to4 I__1310 (
            .O(N__7682),
            .I(N__7679));
    Odrv12 I__1309 (
            .O(N__7679),
            .I(\uu2.mem0.g0_i_a2_4 ));
    InMux I__1308 (
            .O(N__7676),
            .I(N__7673));
    LocalMux I__1307 (
            .O(N__7673),
            .I(\uu2.mem0.N_8_tz_0_0_1 ));
    CascadeMux I__1306 (
            .O(N__7670),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_17_cascade_ ));
    InMux I__1305 (
            .O(N__7667),
            .I(N__7664));
    LocalMux I__1304 (
            .O(N__7664),
            .I(N__7661));
    Odrv4 I__1303 (
            .O(N__7661),
            .I(\uu2.mem0.w_data_5 ));
    InMux I__1302 (
            .O(N__7658),
            .I(N__7652));
    InMux I__1301 (
            .O(N__7657),
            .I(N__7652));
    LocalMux I__1300 (
            .O(N__7652),
            .I(\uu2.Z_decfrac105_7_3 ));
    CascadeMux I__1299 (
            .O(N__7649),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_ ));
    InMux I__1298 (
            .O(N__7646),
            .I(N__7643));
    LocalMux I__1297 (
            .O(N__7643),
            .I(N__7640));
    Span4Mux_h I__1296 (
            .O(N__7640),
            .I(N__7637));
    Odrv4 I__1295 (
            .O(N__7637),
            .I(\uu2.mem0.w_data_0 ));
    InMux I__1294 (
            .O(N__7634),
            .I(N__7631));
    LocalMux I__1293 (
            .O(N__7631),
            .I(N__7628));
    Span4Mux_v I__1292 (
            .O(N__7628),
            .I(N__7625));
    Odrv4 I__1291 (
            .O(N__7625),
            .I(\uu2.mem0.w_data_2 ));
    CascadeMux I__1290 (
            .O(N__7622),
            .I(N__7619));
    InMux I__1289 (
            .O(N__7619),
            .I(N__7616));
    LocalMux I__1288 (
            .O(N__7616),
            .I(\uu2.un1_w_user_cr_0_0 ));
    IoInMux I__1287 (
            .O(N__7613),
            .I(N__7610));
    LocalMux I__1286 (
            .O(N__7610),
            .I(N__7606));
    InMux I__1285 (
            .O(N__7609),
            .I(N__7603));
    Span12Mux_s5_v I__1284 (
            .O(N__7606),
            .I(N__7598));
    LocalMux I__1283 (
            .O(N__7603),
            .I(N__7598));
    Odrv12 I__1282 (
            .O(N__7598),
            .I(latticehx1k_pll_inst_PLLOUTCORE_i));
    CascadeMux I__1281 (
            .O(N__7595),
            .I(\uu2.un1_w_user_cr_0_0_cascade_ ));
    SRMux I__1280 (
            .O(N__7592),
            .I(N__7589));
    LocalMux I__1279 (
            .O(N__7589),
            .I(N__7585));
    CEMux I__1278 (
            .O(N__7588),
            .I(N__7582));
    Span4Mux_v I__1277 (
            .O(N__7585),
            .I(N__7579));
    LocalMux I__1276 (
            .O(N__7582),
            .I(N__7576));
    Span4Mux_h I__1275 (
            .O(N__7579),
            .I(N__7571));
    Span4Mux_v I__1274 (
            .O(N__7576),
            .I(N__7571));
    Span4Mux_s2_h I__1273 (
            .O(N__7571),
            .I(N__7568));
    Odrv4 I__1272 (
            .O(N__7568),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    InMux I__1271 (
            .O(N__7565),
            .I(N__7562));
    LocalMux I__1270 (
            .O(N__7562),
            .I(\resetGen.un3_reset_count_i_a3Z0Z_7 ));
    InMux I__1269 (
            .O(N__7559),
            .I(N__7552));
    InMux I__1268 (
            .O(N__7558),
            .I(N__7552));
    InMux I__1267 (
            .O(N__7557),
            .I(N__7549));
    LocalMux I__1266 (
            .O(N__7552),
            .I(N__7546));
    LocalMux I__1265 (
            .O(N__7549),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    Odrv4 I__1264 (
            .O(N__7546),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    CascadeMux I__1263 (
            .O(N__7541),
            .I(N_87_cascade_));
    InMux I__1262 (
            .O(N__7538),
            .I(N__7534));
    InMux I__1261 (
            .O(N__7537),
            .I(N__7531));
    LocalMux I__1260 (
            .O(N__7534),
            .I(N__7528));
    LocalMux I__1259 (
            .O(N__7531),
            .I(N__7523));
    Span4Mux_v I__1258 (
            .O(N__7528),
            .I(N__7523));
    Odrv4 I__1257 (
            .O(N__7523),
            .I(\buart.Z_rx.N_91 ));
    CascadeMux I__1256 (
            .O(N__7520),
            .I(\buart.Z_rx.N_91_cascade_ ));
    InMux I__1255 (
            .O(N__7517),
            .I(N__7514));
    LocalMux I__1254 (
            .O(N__7514),
            .I(N__7508));
    InMux I__1253 (
            .O(N__7513),
            .I(N__7505));
    InMux I__1252 (
            .O(N__7512),
            .I(N__7500));
    InMux I__1251 (
            .O(N__7511),
            .I(N__7500));
    Odrv4 I__1250 (
            .O(N__7508),
            .I(\buart.Z_rx.N_29_0_i_2 ));
    LocalMux I__1249 (
            .O(N__7505),
            .I(\buart.Z_rx.N_29_0_i_2 ));
    LocalMux I__1248 (
            .O(N__7500),
            .I(\buart.Z_rx.N_29_0_i_2 ));
    InMux I__1247 (
            .O(N__7493),
            .I(N__7490));
    LocalMux I__1246 (
            .O(N__7490),
            .I(N__7487));
    Span4Mux_h I__1245 (
            .O(N__7487),
            .I(N__7484));
    Odrv4 I__1244 (
            .O(N__7484),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    CascadeMux I__1243 (
            .O(N__7481),
            .I(\buart.Z_rx.N_29_0_i_2_cascade_ ));
    CascadeMux I__1242 (
            .O(N__7478),
            .I(N__7475));
    InMux I__1241 (
            .O(N__7475),
            .I(N__7471));
    InMux I__1240 (
            .O(N__7474),
            .I(N__7465));
    LocalMux I__1239 (
            .O(N__7471),
            .I(N__7462));
    InMux I__1238 (
            .O(N__7470),
            .I(N__7455));
    InMux I__1237 (
            .O(N__7469),
            .I(N__7455));
    InMux I__1236 (
            .O(N__7468),
            .I(N__7455));
    LocalMux I__1235 (
            .O(N__7465),
            .I(N__7446));
    Span4Mux_h I__1234 (
            .O(N__7462),
            .I(N__7446));
    LocalMux I__1233 (
            .O(N__7455),
            .I(N__7446));
    InMux I__1232 (
            .O(N__7454),
            .I(N__7437));
    InMux I__1231 (
            .O(N__7453),
            .I(N__7437));
    Span4Mux_v I__1230 (
            .O(N__7446),
            .I(N__7434));
    InMux I__1229 (
            .O(N__7445),
            .I(N__7425));
    InMux I__1228 (
            .O(N__7444),
            .I(N__7425));
    InMux I__1227 (
            .O(N__7443),
            .I(N__7425));
    InMux I__1226 (
            .O(N__7442),
            .I(N__7425));
    LocalMux I__1225 (
            .O(N__7437),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__1224 (
            .O(N__7434),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__1223 (
            .O(N__7425),
            .I(\buart.Z_rx.startbit ));
    CascadeMux I__1222 (
            .O(N__7418),
            .I(N__7414));
    InMux I__1221 (
            .O(N__7417),
            .I(N__7411));
    InMux I__1220 (
            .O(N__7414),
            .I(N__7406));
    LocalMux I__1219 (
            .O(N__7411),
            .I(N__7403));
    InMux I__1218 (
            .O(N__7410),
            .I(N__7398));
    InMux I__1217 (
            .O(N__7409),
            .I(N__7398));
    LocalMux I__1216 (
            .O(N__7406),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    Odrv4 I__1215 (
            .O(N__7403),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    LocalMux I__1214 (
            .O(N__7398),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    CEMux I__1213 (
            .O(N__7391),
            .I(N__7387));
    CEMux I__1212 (
            .O(N__7390),
            .I(N__7384));
    LocalMux I__1211 (
            .O(N__7387),
            .I(N__7380));
    LocalMux I__1210 (
            .O(N__7384),
            .I(N__7377));
    CEMux I__1209 (
            .O(N__7383),
            .I(N__7374));
    Span4Mux_v I__1208 (
            .O(N__7380),
            .I(N__7367));
    Span4Mux_v I__1207 (
            .O(N__7377),
            .I(N__7367));
    LocalMux I__1206 (
            .O(N__7374),
            .I(N__7367));
    Span4Mux_v I__1205 (
            .O(N__7367),
            .I(N__7364));
    Sp12to4 I__1204 (
            .O(N__7364),
            .I(N__7361));
    Odrv12 I__1203 (
            .O(N__7361),
            .I(\buart.Z_rx.bitcounte_0_i_2 ));
    CascadeMux I__1202 (
            .O(N__7358),
            .I(\uu2.Z_decfrac105_7_3_cascade_ ));
    InMux I__1201 (
            .O(N__7355),
            .I(N__7352));
    LocalMux I__1200 (
            .O(N__7352),
            .I(N__7349));
    Odrv12 I__1199 (
            .O(N__7349),
            .I(\uu2.mem0.w_data_6 ));
    InMux I__1198 (
            .O(N__7346),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    InMux I__1197 (
            .O(N__7343),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__1196 (
            .O(N__7340),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    CascadeMux I__1195 (
            .O(N__7337),
            .I(N__7334));
    InMux I__1194 (
            .O(N__7334),
            .I(N__7331));
    LocalMux I__1193 (
            .O(N__7331),
            .I(N__7328));
    Odrv4 I__1192 (
            .O(N__7328),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    CascadeMux I__1191 (
            .O(N__7325),
            .I(N__7322));
    InMux I__1190 (
            .O(N__7322),
            .I(N__7319));
    LocalMux I__1189 (
            .O(N__7319),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__1188 (
            .O(N__7316),
            .I(N__7313));
    LocalMux I__1187 (
            .O(N__7313),
            .I(N__7310));
    Span4Mux_h I__1186 (
            .O(N__7310),
            .I(N__7307));
    Odrv4 I__1185 (
            .O(N__7307),
            .I(\uu2.mem0.w_data_7 ));
    InMux I__1184 (
            .O(N__7304),
            .I(N__7301));
    LocalMux I__1183 (
            .O(N__7301),
            .I(N__7297));
    CascadeMux I__1182 (
            .O(N__7300),
            .I(N__7292));
    Span4Mux_v I__1181 (
            .O(N__7297),
            .I(N__7289));
    InMux I__1180 (
            .O(N__7296),
            .I(N__7282));
    InMux I__1179 (
            .O(N__7295),
            .I(N__7282));
    InMux I__1178 (
            .O(N__7292),
            .I(N__7282));
    Odrv4 I__1177 (
            .O(N__7289),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__1176 (
            .O(N__7282),
            .I(\buart.Z_rx.ser_clk ));
    CascadeMux I__1175 (
            .O(N__7277),
            .I(\buart.Z_rx.N_103_cascade_ ));
    InMux I__1174 (
            .O(N__7274),
            .I(N__7271));
    LocalMux I__1173 (
            .O(N__7271),
            .I(N__7268));
    Span4Mux_v I__1172 (
            .O(N__7268),
            .I(N__7265));
    Odrv4 I__1171 (
            .O(N__7265),
            .I(\uu2.r_data_wire_7 ));
    InMux I__1170 (
            .O(N__7262),
            .I(N__7259));
    LocalMux I__1169 (
            .O(N__7259),
            .I(N__7256));
    Odrv4 I__1168 (
            .O(N__7256),
            .I(vbuf_tx_data_7));
    CEMux I__1167 (
            .O(N__7253),
            .I(N__7250));
    LocalMux I__1166 (
            .O(N__7250),
            .I(N__7247));
    Span4Mux_v I__1165 (
            .O(N__7247),
            .I(N__7243));
    CEMux I__1164 (
            .O(N__7246),
            .I(N__7240));
    Odrv4 I__1163 (
            .O(N__7243),
            .I(\uu2.vbuf_tx_data_rdy_0 ));
    LocalMux I__1162 (
            .O(N__7240),
            .I(\uu2.vbuf_tx_data_rdy_0 ));
    InMux I__1161 (
            .O(N__7235),
            .I(N__7232));
    LocalMux I__1160 (
            .O(N__7232),
            .I(vbuf_tx_data_3));
    InMux I__1159 (
            .O(N__7229),
            .I(N__7226));
    LocalMux I__1158 (
            .O(N__7226),
            .I(vbuf_tx_data_4));
    InMux I__1157 (
            .O(N__7223),
            .I(N__7220));
    LocalMux I__1156 (
            .O(N__7220),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    CascadeMux I__1155 (
            .O(N__7217),
            .I(N__7214));
    InMux I__1154 (
            .O(N__7214),
            .I(N__7211));
    LocalMux I__1153 (
            .O(N__7211),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__1152 (
            .O(N__7208),
            .I(N__7205));
    LocalMux I__1151 (
            .O(N__7205),
            .I(vbuf_tx_data_2));
    CascadeMux I__1150 (
            .O(N__7202),
            .I(N__7199));
    InMux I__1149 (
            .O(N__7199),
            .I(N__7196));
    LocalMux I__1148 (
            .O(N__7196),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__1147 (
            .O(N__7193),
            .I(N__7190));
    LocalMux I__1146 (
            .O(N__7190),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__1145 (
            .O(N__7187),
            .I(N__7184));
    LocalMux I__1144 (
            .O(N__7184),
            .I(N__7181));
    IoSpan4Mux I__1143 (
            .O(N__7181),
            .I(N__7178));
    Span4Mux_s3_h I__1142 (
            .O(N__7178),
            .I(N__7175));
    Odrv4 I__1141 (
            .O(N__7175),
            .I(o_serial_data_c));
    InMux I__1140 (
            .O(N__7172),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    CascadeMux I__1139 (
            .O(N__7169),
            .I(\buart.Z_rx.ser_clk_cascade_ ));
    InMux I__1138 (
            .O(N__7166),
            .I(N__7163));
    LocalMux I__1137 (
            .O(N__7163),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    CascadeMux I__1136 (
            .O(N__7160),
            .I(N__7157));
    InMux I__1135 (
            .O(N__7157),
            .I(N__7152));
    InMux I__1134 (
            .O(N__7156),
            .I(N__7147));
    InMux I__1133 (
            .O(N__7155),
            .I(N__7147));
    LocalMux I__1132 (
            .O(N__7152),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__1131 (
            .O(N__7147),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    InMux I__1130 (
            .O(N__7142),
            .I(N__7139));
    LocalMux I__1129 (
            .O(N__7139),
            .I(N__7136));
    Span4Mux_h I__1128 (
            .O(N__7136),
            .I(N__7133));
    Span4Mux_v I__1127 (
            .O(N__7133),
            .I(N__7130));
    Odrv4 I__1126 (
            .O(N__7130),
            .I(\uu2.r_data_wire_0 ));
    InMux I__1125 (
            .O(N__7127),
            .I(N__7124));
    LocalMux I__1124 (
            .O(N__7124),
            .I(N__7121));
    Span4Mux_h I__1123 (
            .O(N__7121),
            .I(N__7118));
    Span4Mux_v I__1122 (
            .O(N__7118),
            .I(N__7115));
    Odrv4 I__1121 (
            .O(N__7115),
            .I(\uu2.r_data_wire_1 ));
    InMux I__1120 (
            .O(N__7112),
            .I(N__7109));
    LocalMux I__1119 (
            .O(N__7109),
            .I(N__7106));
    Span4Mux_v I__1118 (
            .O(N__7106),
            .I(N__7103));
    Span4Mux_v I__1117 (
            .O(N__7103),
            .I(N__7100));
    Odrv4 I__1116 (
            .O(N__7100),
            .I(\uu2.r_data_wire_2 ));
    InMux I__1115 (
            .O(N__7097),
            .I(N__7094));
    LocalMux I__1114 (
            .O(N__7094),
            .I(N__7091));
    Span12Mux_s9_v I__1113 (
            .O(N__7091),
            .I(N__7088));
    Odrv12 I__1112 (
            .O(N__7088),
            .I(\uu2.r_data_wire_3 ));
    InMux I__1111 (
            .O(N__7085),
            .I(N__7082));
    LocalMux I__1110 (
            .O(N__7082),
            .I(N__7079));
    Span4Mux_v I__1109 (
            .O(N__7079),
            .I(N__7076));
    Odrv4 I__1108 (
            .O(N__7076),
            .I(\uu2.r_data_wire_4 ));
    InMux I__1107 (
            .O(N__7073),
            .I(N__7070));
    LocalMux I__1106 (
            .O(N__7070),
            .I(N__7067));
    Span4Mux_h I__1105 (
            .O(N__7067),
            .I(N__7064));
    Span4Mux_v I__1104 (
            .O(N__7064),
            .I(N__7061));
    Odrv4 I__1103 (
            .O(N__7061),
            .I(\uu2.r_data_wire_5 ));
    InMux I__1102 (
            .O(N__7058),
            .I(N__7055));
    LocalMux I__1101 (
            .O(N__7055),
            .I(N__7052));
    Odrv4 I__1100 (
            .O(N__7052),
            .I(vbuf_tx_data_5));
    InMux I__1099 (
            .O(N__7049),
            .I(N__7046));
    LocalMux I__1098 (
            .O(N__7046),
            .I(N__7043));
    Span12Mux_s9_h I__1097 (
            .O(N__7043),
            .I(N__7040));
    Odrv12 I__1096 (
            .O(N__7040),
            .I(\uu2.r_data_wire_6 ));
    InMux I__1095 (
            .O(N__7037),
            .I(N__7034));
    LocalMux I__1094 (
            .O(N__7034),
            .I(vbuf_tx_data_6));
    InMux I__1093 (
            .O(N__7031),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    InMux I__1092 (
            .O(N__7028),
            .I(N__7025));
    LocalMux I__1091 (
            .O(N__7025),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    CascadeMux I__1090 (
            .O(N__7022),
            .I(N__7019));
    InMux I__1089 (
            .O(N__7019),
            .I(N__7016));
    LocalMux I__1088 (
            .O(N__7016),
            .I(N__7013));
    Span4Mux_h I__1087 (
            .O(N__7013),
            .I(N__7010));
    Odrv4 I__1086 (
            .O(N__7010),
            .I(\uu2.mem0.g0_0_a3_0 ));
    CascadeMux I__1085 (
            .O(N__7007),
            .I(\buart.Z_rx.startbit_cascade_ ));
    InMux I__1084 (
            .O(N__7004),
            .I(N__6998));
    InMux I__1083 (
            .O(N__7003),
            .I(N__6998));
    LocalMux I__1082 (
            .O(N__6998),
            .I(N__6995));
    Odrv4 I__1081 (
            .O(N__6995),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    InMux I__1080 (
            .O(N__6992),
            .I(N__6988));
    InMux I__1079 (
            .O(N__6991),
            .I(N__6985));
    LocalMux I__1078 (
            .O(N__6988),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__1077 (
            .O(N__6985),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    CascadeMux I__1076 (
            .O(N__6980),
            .I(N__6977));
    InMux I__1075 (
            .O(N__6977),
            .I(N__6970));
    InMux I__1074 (
            .O(N__6976),
            .I(N__6970));
    InMux I__1073 (
            .O(N__6975),
            .I(N__6967));
    LocalMux I__1072 (
            .O(N__6970),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__1071 (
            .O(N__6967),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__1070 (
            .O(N__6962),
            .I(N__6958));
    CascadeMux I__1069 (
            .O(N__6961),
            .I(N__6955));
    InMux I__1068 (
            .O(N__6958),
            .I(N__6952));
    InMux I__1067 (
            .O(N__6955),
            .I(N__6949));
    LocalMux I__1066 (
            .O(N__6952),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    LocalMux I__1065 (
            .O(N__6949),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    InMux I__1064 (
            .O(N__6944),
            .I(N__6939));
    InMux I__1063 (
            .O(N__6943),
            .I(N__6934));
    InMux I__1062 (
            .O(N__6942),
            .I(N__6934));
    LocalMux I__1061 (
            .O(N__6939),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1060 (
            .O(N__6934),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__1059 (
            .O(N__6929),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ));
    CascadeMux I__1058 (
            .O(N__6926),
            .I(N__6920));
    InMux I__1057 (
            .O(N__6925),
            .I(N__6913));
    InMux I__1056 (
            .O(N__6924),
            .I(N__6913));
    InMux I__1055 (
            .O(N__6923),
            .I(N__6913));
    InMux I__1054 (
            .O(N__6920),
            .I(N__6910));
    LocalMux I__1053 (
            .O(N__6913),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1052 (
            .O(N__6910),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__1051 (
            .O(N__6905),
            .I(N__6902));
    LocalMux I__1050 (
            .O(N__6902),
            .I(\uu2.mem0.g0_i_5 ));
    InMux I__1049 (
            .O(N__6899),
            .I(N__6896));
    LocalMux I__1048 (
            .O(N__6896),
            .I(\uu2.mem0.g0_i_6_1_0 ));
    CascadeMux I__1047 (
            .O(N__6893),
            .I(\uu2.mem0.N_19_cascade_ ));
    InMux I__1046 (
            .O(N__6890),
            .I(N__6887));
    LocalMux I__1045 (
            .O(N__6887),
            .I(\uu2.mem0.g0_i_6 ));
    InMux I__1044 (
            .O(N__6884),
            .I(N__6881));
    LocalMux I__1043 (
            .O(N__6881),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_53 ));
    InMux I__1042 (
            .O(N__6878),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__1041 (
            .O(N__6875),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__1040 (
            .O(N__6872),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    CascadeMux I__1039 (
            .O(N__6869),
            .I(\uu2.mem0.g2_1_0_0_cascade_ ));
    InMux I__1038 (
            .O(N__6866),
            .I(N__6863));
    LocalMux I__1037 (
            .O(N__6863),
            .I(\uu2.mem0.g0_2_1 ));
    CascadeMux I__1036 (
            .O(N__6860),
            .I(\uu2.mem0.g0_i_a2_3_cascade_ ));
    InMux I__1035 (
            .O(N__6857),
            .I(N__6854));
    LocalMux I__1034 (
            .O(N__6854),
            .I(\uu2.mem0.w_data_displaying_2_0_0 ));
    InMux I__1033 (
            .O(N__6851),
            .I(N__6848));
    LocalMux I__1032 (
            .O(N__6848),
            .I(\uu2.mem0.g1_0_5 ));
    InMux I__1031 (
            .O(N__6845),
            .I(N__6842));
    LocalMux I__1030 (
            .O(N__6842),
            .I(\uu2.mem0.N_10_0_0 ));
    InMux I__1029 (
            .O(N__6839),
            .I(N__6836));
    LocalMux I__1028 (
            .O(N__6836),
            .I(N__6833));
    Odrv4 I__1027 (
            .O(N__6833),
            .I(\uu2.mem0.g1_2 ));
    CascadeMux I__1026 (
            .O(N__6830),
            .I(N__6827));
    InMux I__1025 (
            .O(N__6827),
            .I(N__6824));
    LocalMux I__1024 (
            .O(N__6824),
            .I(\uu2.mem0.g1_1_sx ));
    InMux I__1023 (
            .O(N__6821),
            .I(N__6818));
    LocalMux I__1022 (
            .O(N__6818),
            .I(N__6815));
    Odrv4 I__1021 (
            .O(N__6815),
            .I(\uu2.mem0.g1_0 ));
    CascadeMux I__1020 (
            .O(N__6812),
            .I(\resetGen.N_104_cascade_ ));
    InMux I__1019 (
            .O(N__6809),
            .I(N__6806));
    LocalMux I__1018 (
            .O(N__6806),
            .I(\resetGen.N_84 ));
    InMux I__1017 (
            .O(N__6803),
            .I(N__6791));
    InMux I__1016 (
            .O(N__6802),
            .I(N__6791));
    InMux I__1015 (
            .O(N__6801),
            .I(N__6791));
    InMux I__1014 (
            .O(N__6800),
            .I(N__6791));
    LocalMux I__1013 (
            .O(N__6791),
            .I(\resetGen.reset_countZ0Z_0 ));
    InMux I__1012 (
            .O(N__6788),
            .I(N__6779));
    InMux I__1011 (
            .O(N__6787),
            .I(N__6779));
    InMux I__1010 (
            .O(N__6786),
            .I(N__6779));
    LocalMux I__1009 (
            .O(N__6779),
            .I(\resetGen.reset_countZ0Z_1 ));
    CascadeMux I__1008 (
            .O(N__6776),
            .I(N__6773));
    InMux I__1007 (
            .O(N__6773),
            .I(N__6769));
    InMux I__1006 (
            .O(N__6772),
            .I(N__6766));
    LocalMux I__1005 (
            .O(N__6769),
            .I(\resetGen.reset_countZ0Z_2 ));
    LocalMux I__1004 (
            .O(N__6766),
            .I(\resetGen.reset_countZ0Z_2 ));
    InMux I__1003 (
            .O(N__6761),
            .I(N__6758));
    LocalMux I__1002 (
            .O(N__6758),
            .I(\resetGen.N_86 ));
    InMux I__1001 (
            .O(N__6755),
            .I(N__6743));
    InMux I__1000 (
            .O(N__6754),
            .I(N__6743));
    InMux I__999 (
            .O(N__6753),
            .I(N__6743));
    InMux I__998 (
            .O(N__6752),
            .I(N__6743));
    LocalMux I__997 (
            .O(N__6743),
            .I(\resetGen.N_104 ));
    InMux I__996 (
            .O(N__6740),
            .I(N__6734));
    InMux I__995 (
            .O(N__6739),
            .I(N__6734));
    LocalMux I__994 (
            .O(N__6734),
            .I(\resetGen.reset_countZ0Z_3 ));
    CascadeMux I__993 (
            .O(N__6731),
            .I(\resetGen.N_86_cascade_ ));
    InMux I__992 (
            .O(N__6728),
            .I(N__6724));
    CascadeMux I__991 (
            .O(N__6727),
            .I(N__6720));
    LocalMux I__990 (
            .O(N__6724),
            .I(N__6714));
    InMux I__989 (
            .O(N__6723),
            .I(N__6710));
    InMux I__988 (
            .O(N__6720),
            .I(N__6701));
    InMux I__987 (
            .O(N__6719),
            .I(N__6701));
    InMux I__986 (
            .O(N__6718),
            .I(N__6701));
    InMux I__985 (
            .O(N__6717),
            .I(N__6701));
    Span4Mux_h I__984 (
            .O(N__6714),
            .I(N__6698));
    InMux I__983 (
            .O(N__6713),
            .I(N__6695));
    LocalMux I__982 (
            .O(N__6710),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__981 (
            .O(N__6701),
            .I(\resetGen.reset_countZ0Z_4 ));
    Odrv4 I__980 (
            .O(N__6698),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__979 (
            .O(N__6695),
            .I(\resetGen.reset_countZ0Z_4 ));
    InMux I__978 (
            .O(N__6686),
            .I(N__6683));
    LocalMux I__977 (
            .O(N__6683),
            .I(\Lab_UT.secuu0.un4_l_count_12 ));
    CascadeMux I__976 (
            .O(N__6680),
            .I(N__6677));
    InMux I__975 (
            .O(N__6677),
            .I(N__6674));
    LocalMux I__974 (
            .O(N__6674),
            .I(\Lab_UT.secuu0.un87_ci ));
    CascadeMux I__973 (
            .O(N__6671),
            .I(\Lab_UT.secuu0.un87_ci_cascade_ ));
    InMux I__972 (
            .O(N__6668),
            .I(N__6661));
    InMux I__971 (
            .O(N__6667),
            .I(N__6661));
    InMux I__970 (
            .O(N__6666),
            .I(N__6658));
    LocalMux I__969 (
            .O(N__6661),
            .I(\Lab_UT.secuu0.l_countZ0Z_3 ));
    LocalMux I__968 (
            .O(N__6658),
            .I(\Lab_UT.secuu0.l_countZ0Z_3 ));
    InMux I__967 (
            .O(N__6653),
            .I(N__6643));
    InMux I__966 (
            .O(N__6652),
            .I(N__6643));
    InMux I__965 (
            .O(N__6651),
            .I(N__6643));
    InMux I__964 (
            .O(N__6650),
            .I(N__6640));
    LocalMux I__963 (
            .O(N__6643),
            .I(\Lab_UT.secuu0.l_countZ0Z_2 ));
    LocalMux I__962 (
            .O(N__6640),
            .I(\Lab_UT.secuu0.l_countZ0Z_2 ));
    CascadeMux I__961 (
            .O(N__6635),
            .I(N__6629));
    InMux I__960 (
            .O(N__6634),
            .I(N__6625));
    InMux I__959 (
            .O(N__6633),
            .I(N__6618));
    InMux I__958 (
            .O(N__6632),
            .I(N__6618));
    InMux I__957 (
            .O(N__6629),
            .I(N__6618));
    InMux I__956 (
            .O(N__6628),
            .I(N__6615));
    LocalMux I__955 (
            .O(N__6625),
            .I(\Lab_UT.secuu0.l_countZ0Z_0 ));
    LocalMux I__954 (
            .O(N__6618),
            .I(\Lab_UT.secuu0.l_countZ0Z_0 ));
    LocalMux I__953 (
            .O(N__6615),
            .I(\Lab_UT.secuu0.l_countZ0Z_0 ));
    InMux I__952 (
            .O(N__6608),
            .I(N__6602));
    InMux I__951 (
            .O(N__6607),
            .I(N__6595));
    InMux I__950 (
            .O(N__6606),
            .I(N__6595));
    InMux I__949 (
            .O(N__6605),
            .I(N__6595));
    LocalMux I__948 (
            .O(N__6602),
            .I(N__6592));
    LocalMux I__947 (
            .O(N__6595),
            .I(\Lab_UT.secuu0.l_countZ0Z_1 ));
    Odrv4 I__946 (
            .O(N__6592),
            .I(\Lab_UT.secuu0.l_countZ0Z_1 ));
    CascadeMux I__945 (
            .O(N__6587),
            .I(\Lab_UT.secuu0.un109_ci_cascade_ ));
    CascadeMux I__944 (
            .O(N__6584),
            .I(N__6578));
    CascadeMux I__943 (
            .O(N__6583),
            .I(N__6569));
    InMux I__942 (
            .O(N__6582),
            .I(N__6565));
    InMux I__941 (
            .O(N__6581),
            .I(N__6562));
    InMux I__940 (
            .O(N__6578),
            .I(N__6557));
    InMux I__939 (
            .O(N__6577),
            .I(N__6557));
    InMux I__938 (
            .O(N__6576),
            .I(N__6546));
    InMux I__937 (
            .O(N__6575),
            .I(N__6546));
    InMux I__936 (
            .O(N__6574),
            .I(N__6546));
    InMux I__935 (
            .O(N__6573),
            .I(N__6546));
    InMux I__934 (
            .O(N__6572),
            .I(N__6546));
    InMux I__933 (
            .O(N__6569),
            .I(N__6541));
    InMux I__932 (
            .O(N__6568),
            .I(N__6541));
    LocalMux I__931 (
            .O(N__6565),
            .I(\Lab_UT.secuu0.un153_ci ));
    LocalMux I__930 (
            .O(N__6562),
            .I(\Lab_UT.secuu0.un153_ci ));
    LocalMux I__929 (
            .O(N__6557),
            .I(\Lab_UT.secuu0.un153_ci ));
    LocalMux I__928 (
            .O(N__6546),
            .I(\Lab_UT.secuu0.un153_ci ));
    LocalMux I__927 (
            .O(N__6541),
            .I(\Lab_UT.secuu0.un153_ci ));
    InMux I__926 (
            .O(N__6530),
            .I(N__6524));
    InMux I__925 (
            .O(N__6529),
            .I(N__6524));
    LocalMux I__924 (
            .O(N__6524),
            .I(N__6521));
    Odrv4 I__923 (
            .O(N__6521),
            .I(\Lab_UT.secuu0.un131_ci_3 ));
    InMux I__922 (
            .O(N__6518),
            .I(N__6514));
    InMux I__921 (
            .O(N__6517),
            .I(N__6509));
    LocalMux I__920 (
            .O(N__6514),
            .I(N__6506));
    InMux I__919 (
            .O(N__6513),
            .I(N__6501));
    InMux I__918 (
            .O(N__6512),
            .I(N__6501));
    LocalMux I__917 (
            .O(N__6509),
            .I(N__6498));
    Odrv4 I__916 (
            .O(N__6506),
            .I(\Lab_UT.secuu0.l_countZ0Z_6 ));
    LocalMux I__915 (
            .O(N__6501),
            .I(\Lab_UT.secuu0.l_countZ0Z_6 ));
    Odrv4 I__914 (
            .O(N__6498),
            .I(\Lab_UT.secuu0.l_countZ0Z_6 ));
    CascadeMux I__913 (
            .O(N__6491),
            .I(N__6488));
    InMux I__912 (
            .O(N__6488),
            .I(N__6477));
    InMux I__911 (
            .O(N__6487),
            .I(N__6477));
    InMux I__910 (
            .O(N__6486),
            .I(N__6472));
    InMux I__909 (
            .O(N__6485),
            .I(N__6472));
    InMux I__908 (
            .O(N__6484),
            .I(N__6465));
    InMux I__907 (
            .O(N__6483),
            .I(N__6465));
    InMux I__906 (
            .O(N__6482),
            .I(N__6465));
    LocalMux I__905 (
            .O(N__6477),
            .I(N__6453));
    LocalMux I__904 (
            .O(N__6472),
            .I(N__6453));
    LocalMux I__903 (
            .O(N__6465),
            .I(N__6453));
    InMux I__902 (
            .O(N__6464),
            .I(N__6450));
    InMux I__901 (
            .O(N__6463),
            .I(N__6441));
    InMux I__900 (
            .O(N__6462),
            .I(N__6441));
    InMux I__899 (
            .O(N__6461),
            .I(N__6441));
    InMux I__898 (
            .O(N__6460),
            .I(N__6441));
    Odrv4 I__897 (
            .O(N__6453),
            .I(\Lab_UT.secuu0.un4_l_count_0 ));
    LocalMux I__896 (
            .O(N__6450),
            .I(\Lab_UT.secuu0.un4_l_count_0 ));
    LocalMux I__895 (
            .O(N__6441),
            .I(\Lab_UT.secuu0.un4_l_count_0 ));
    InMux I__894 (
            .O(N__6434),
            .I(N__6431));
    LocalMux I__893 (
            .O(N__6431),
            .I(N__6428));
    Odrv12 I__892 (
            .O(N__6428),
            .I(\Lab_UT.secuu0.un142_ci_0 ));
    InMux I__891 (
            .O(N__6425),
            .I(N__6422));
    LocalMux I__890 (
            .O(N__6422),
            .I(N__6418));
    CascadeMux I__889 (
            .O(N__6421),
            .I(N__6413));
    Span4Mux_h I__888 (
            .O(N__6418),
            .I(N__6410));
    InMux I__887 (
            .O(N__6417),
            .I(N__6407));
    InMux I__886 (
            .O(N__6416),
            .I(N__6402));
    InMux I__885 (
            .O(N__6413),
            .I(N__6402));
    Odrv4 I__884 (
            .O(N__6410),
            .I(\Lab_UT.secuu0.un109_ci ));
    LocalMux I__883 (
            .O(N__6407),
            .I(\Lab_UT.secuu0.un109_ci ));
    LocalMux I__882 (
            .O(N__6402),
            .I(\Lab_UT.secuu0.un109_ci ));
    CascadeMux I__881 (
            .O(N__6395),
            .I(N__6392));
    InMux I__880 (
            .O(N__6392),
            .I(N__6387));
    InMux I__879 (
            .O(N__6391),
            .I(N__6384));
    InMux I__878 (
            .O(N__6390),
            .I(N__6381));
    LocalMux I__877 (
            .O(N__6387),
            .I(\Lab_UT.secuu0.l_countZ0Z_7 ));
    LocalMux I__876 (
            .O(N__6384),
            .I(\Lab_UT.secuu0.l_countZ0Z_7 ));
    LocalMux I__875 (
            .O(N__6381),
            .I(\Lab_UT.secuu0.l_countZ0Z_7 ));
    CEMux I__874 (
            .O(N__6374),
            .I(N__6359));
    CEMux I__873 (
            .O(N__6373),
            .I(N__6359));
    CEMux I__872 (
            .O(N__6372),
            .I(N__6359));
    CEMux I__871 (
            .O(N__6371),
            .I(N__6359));
    CEMux I__870 (
            .O(N__6370),
            .I(N__6359));
    GlobalMux I__869 (
            .O(N__6359),
            .I(N__6356));
    gio2CtrlBuf I__868 (
            .O(N__6356),
            .I(\Lab_UT.secuu0.un11_l_count_i_g ));
    InMux I__867 (
            .O(N__6353),
            .I(N__6350));
    LocalMux I__866 (
            .O(N__6350),
            .I(\Lab_UT.secuu0.un4_l_count_13 ));
    CascadeMux I__865 (
            .O(N__6347),
            .I(\Lab_UT.secuu0.un4_l_count_16_cascade_ ));
    InMux I__864 (
            .O(N__6344),
            .I(N__6341));
    LocalMux I__863 (
            .O(N__6341),
            .I(N__6338));
    Odrv4 I__862 (
            .O(N__6338),
            .I(\Lab_UT.secuu0.un4_l_count_18 ));
    InMux I__861 (
            .O(N__6335),
            .I(N__6332));
    LocalMux I__860 (
            .O(N__6332),
            .I(\Lab_UT.secuu0.delay_lineZ0Z_1 ));
    CascadeMux I__859 (
            .O(N__6329),
            .I(\Lab_UT.secuu0.un4_l_count_0_cascade_ ));
    InMux I__858 (
            .O(N__6326),
            .I(N__6322));
    InMux I__857 (
            .O(N__6325),
            .I(N__6319));
    LocalMux I__856 (
            .O(N__6322),
            .I(\Lab_UT.secuu0.delay_lineZ0Z_0 ));
    LocalMux I__855 (
            .O(N__6319),
            .I(\Lab_UT.secuu0.delay_lineZ0Z_0 ));
    IoInMux I__854 (
            .O(N__6314),
            .I(N__6311));
    LocalMux I__853 (
            .O(N__6311),
            .I(N__6308));
    IoSpan4Mux I__852 (
            .O(N__6308),
            .I(N__6305));
    Span4Mux_s0_h I__851 (
            .O(N__6305),
            .I(N__6302));
    Span4Mux_h I__850 (
            .O(N__6302),
            .I(N__6299));
    Odrv4 I__849 (
            .O(N__6299),
            .I(\Lab_UT.secuu0.un11_l_count_i ));
    CascadeMux I__848 (
            .O(N__6296),
            .I(N__6293));
    InMux I__847 (
            .O(N__6293),
            .I(N__6290));
    LocalMux I__846 (
            .O(N__6290),
            .I(\Lab_UT.secuu0.un186_ci_0 ));
    InMux I__845 (
            .O(N__6287),
            .I(N__6282));
    InMux I__844 (
            .O(N__6286),
            .I(N__6279));
    InMux I__843 (
            .O(N__6285),
            .I(N__6276));
    LocalMux I__842 (
            .O(N__6282),
            .I(\Lab_UT.secuu0.l_countZ0Z_11 ));
    LocalMux I__841 (
            .O(N__6279),
            .I(\Lab_UT.secuu0.l_countZ0Z_11 ));
    LocalMux I__840 (
            .O(N__6276),
            .I(\Lab_UT.secuu0.l_countZ0Z_11 ));
    CascadeMux I__839 (
            .O(N__6269),
            .I(N__6264));
    InMux I__838 (
            .O(N__6268),
            .I(N__6257));
    InMux I__837 (
            .O(N__6267),
            .I(N__6257));
    InMux I__836 (
            .O(N__6264),
            .I(N__6257));
    LocalMux I__835 (
            .O(N__6257),
            .I(\Lab_UT.secuu0.un241_ci_2 ));
    InMux I__834 (
            .O(N__6254),
            .I(N__6248));
    InMux I__833 (
            .O(N__6253),
            .I(N__6241));
    InMux I__832 (
            .O(N__6252),
            .I(N__6241));
    InMux I__831 (
            .O(N__6251),
            .I(N__6241));
    LocalMux I__830 (
            .O(N__6248),
            .I(N__6238));
    LocalMux I__829 (
            .O(N__6241),
            .I(\Lab_UT.secuu0.l_countZ0Z_16 ));
    Odrv4 I__828 (
            .O(N__6238),
            .I(\Lab_UT.secuu0.l_countZ0Z_16 ));
    CascadeMux I__827 (
            .O(N__6233),
            .I(\Lab_UT.secuu0.un263_ci_cascade_ ));
    InMux I__826 (
            .O(N__6230),
            .I(N__6226));
    InMux I__825 (
            .O(N__6229),
            .I(N__6223));
    LocalMux I__824 (
            .O(N__6226),
            .I(\Lab_UT.secuu0.l_countZ0Z_18 ));
    LocalMux I__823 (
            .O(N__6223),
            .I(\Lab_UT.secuu0.l_countZ0Z_18 ));
    CascadeMux I__822 (
            .O(N__6218),
            .I(N__6214));
    CascadeMux I__821 (
            .O(N__6217),
            .I(N__6209));
    InMux I__820 (
            .O(N__6214),
            .I(N__6205));
    InMux I__819 (
            .O(N__6213),
            .I(N__6198));
    InMux I__818 (
            .O(N__6212),
            .I(N__6198));
    InMux I__817 (
            .O(N__6209),
            .I(N__6198));
    InMux I__816 (
            .O(N__6208),
            .I(N__6195));
    LocalMux I__815 (
            .O(N__6205),
            .I(\Lab_UT.secuu0.l_countZ0Z_9 ));
    LocalMux I__814 (
            .O(N__6198),
            .I(\Lab_UT.secuu0.l_countZ0Z_9 ));
    LocalMux I__813 (
            .O(N__6195),
            .I(\Lab_UT.secuu0.l_countZ0Z_9 ));
    CascadeMux I__812 (
            .O(N__6188),
            .I(N__6183));
    InMux I__811 (
            .O(N__6187),
            .I(N__6176));
    InMux I__810 (
            .O(N__6186),
            .I(N__6176));
    InMux I__809 (
            .O(N__6183),
            .I(N__6176));
    LocalMux I__808 (
            .O(N__6176),
            .I(\Lab_UT.secuu0.l_countZ0Z_17 ));
    InMux I__807 (
            .O(N__6173),
            .I(N__6169));
    InMux I__806 (
            .O(N__6172),
            .I(N__6165));
    LocalMux I__805 (
            .O(N__6169),
            .I(N__6162));
    InMux I__804 (
            .O(N__6168),
            .I(N__6159));
    LocalMux I__803 (
            .O(N__6165),
            .I(\uu2.l_countZ0Z_7 ));
    Odrv4 I__802 (
            .O(N__6162),
            .I(\uu2.l_countZ0Z_7 ));
    LocalMux I__801 (
            .O(N__6159),
            .I(\uu2.l_countZ0Z_7 ));
    CascadeMux I__800 (
            .O(N__6152),
            .I(N__6148));
    CascadeMux I__799 (
            .O(N__6151),
            .I(N__6145));
    InMux I__798 (
            .O(N__6148),
            .I(N__6140));
    InMux I__797 (
            .O(N__6145),
            .I(N__6140));
    LocalMux I__796 (
            .O(N__6140),
            .I(\uu2.vbuf_count.un372_ci_8_1 ));
    CascadeMux I__795 (
            .O(N__6137),
            .I(N__6131));
    InMux I__794 (
            .O(N__6136),
            .I(N__6124));
    InMux I__793 (
            .O(N__6135),
            .I(N__6124));
    InMux I__792 (
            .O(N__6134),
            .I(N__6124));
    InMux I__791 (
            .O(N__6131),
            .I(N__6121));
    LocalMux I__790 (
            .O(N__6124),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__789 (
            .O(N__6121),
            .I(\uu2.l_countZ0Z_8 ));
    CascadeMux I__788 (
            .O(N__6116),
            .I(\uu2.vbuf_count.un372_ci_8_1_cascade_ ));
    InMux I__787 (
            .O(N__6113),
            .I(N__6106));
    InMux I__786 (
            .O(N__6112),
            .I(N__6106));
    InMux I__785 (
            .O(N__6111),
            .I(N__6103));
    LocalMux I__784 (
            .O(N__6106),
            .I(\uu2.l_countZ0Z_9 ));
    LocalMux I__783 (
            .O(N__6103),
            .I(\uu2.l_countZ0Z_9 ));
    InMux I__782 (
            .O(N__6098),
            .I(N__6094));
    InMux I__781 (
            .O(N__6097),
            .I(N__6089));
    LocalMux I__780 (
            .O(N__6094),
            .I(N__6086));
    InMux I__779 (
            .O(N__6093),
            .I(N__6081));
    InMux I__778 (
            .O(N__6092),
            .I(N__6081));
    LocalMux I__777 (
            .O(N__6089),
            .I(N__6078));
    Odrv4 I__776 (
            .O(N__6086),
            .I(\uu2.l_countZ0Z_6 ));
    LocalMux I__775 (
            .O(N__6081),
            .I(\uu2.l_countZ0Z_6 ));
    Odrv4 I__774 (
            .O(N__6078),
            .I(\uu2.l_countZ0Z_6 ));
    InMux I__773 (
            .O(N__6071),
            .I(N__6068));
    LocalMux I__772 (
            .O(N__6068),
            .I(N__6061));
    InMux I__771 (
            .O(N__6067),
            .I(N__6054));
    InMux I__770 (
            .O(N__6066),
            .I(N__6054));
    InMux I__769 (
            .O(N__6065),
            .I(N__6054));
    InMux I__768 (
            .O(N__6064),
            .I(N__6051));
    Odrv4 I__767 (
            .O(N__6061),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__766 (
            .O(N__6054),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__765 (
            .O(N__6051),
            .I(\uu2.l_countZ0Z_5 ));
    CascadeMux I__764 (
            .O(N__6044),
            .I(N__6040));
    InMux I__763 (
            .O(N__6043),
            .I(N__6023));
    InMux I__762 (
            .O(N__6040),
            .I(N__6023));
    InMux I__761 (
            .O(N__6039),
            .I(N__6023));
    InMux I__760 (
            .O(N__6038),
            .I(N__6023));
    InMux I__759 (
            .O(N__6037),
            .I(N__6023));
    InMux I__758 (
            .O(N__6036),
            .I(N__6023));
    LocalMux I__757 (
            .O(N__6023),
            .I(N__6020));
    Odrv4 I__756 (
            .O(N__6020),
            .I(\uu2.un306_ci ));
    CascadeMux I__755 (
            .O(N__6017),
            .I(N__6010));
    CascadeMux I__754 (
            .O(N__6016),
            .I(N__6006));
    CascadeMux I__753 (
            .O(N__6015),
            .I(N__6003));
    InMux I__752 (
            .O(N__6014),
            .I(N__6000));
    InMux I__751 (
            .O(N__6013),
            .I(N__5997));
    InMux I__750 (
            .O(N__6010),
            .I(N__5988));
    InMux I__749 (
            .O(N__6009),
            .I(N__5988));
    InMux I__748 (
            .O(N__6006),
            .I(N__5988));
    InMux I__747 (
            .O(N__6003),
            .I(N__5988));
    LocalMux I__746 (
            .O(N__6000),
            .I(N__5983));
    LocalMux I__745 (
            .O(N__5997),
            .I(N__5983));
    LocalMux I__744 (
            .O(N__5988),
            .I(\uu2.l_countZ0Z_4 ));
    Odrv12 I__743 (
            .O(N__5983),
            .I(\uu2.l_countZ0Z_4 ));
    CascadeMux I__742 (
            .O(N__5978),
            .I(N__5972));
    InMux I__741 (
            .O(N__5977),
            .I(N__5965));
    InMux I__740 (
            .O(N__5976),
            .I(N__5965));
    InMux I__739 (
            .O(N__5975),
            .I(N__5965));
    InMux I__738 (
            .O(N__5972),
            .I(N__5962));
    LocalMux I__737 (
            .O(N__5965),
            .I(\Lab_UT.secuu0.l_precountZ0Z_2 ));
    LocalMux I__736 (
            .O(N__5962),
            .I(\Lab_UT.secuu0.l_precountZ0Z_2 ));
    InMux I__735 (
            .O(N__5957),
            .I(N__5944));
    InMux I__734 (
            .O(N__5956),
            .I(N__5944));
    InMux I__733 (
            .O(N__5955),
            .I(N__5944));
    InMux I__732 (
            .O(N__5954),
            .I(N__5944));
    InMux I__731 (
            .O(N__5953),
            .I(N__5941));
    LocalMux I__730 (
            .O(N__5944),
            .I(\Lab_UT.secuu0.l_precountZ0Z_1 ));
    LocalMux I__729 (
            .O(N__5941),
            .I(\Lab_UT.secuu0.l_precountZ0Z_1 ));
    InMux I__728 (
            .O(N__5936),
            .I(N__5932));
    InMux I__727 (
            .O(N__5935),
            .I(N__5928));
    LocalMux I__726 (
            .O(N__5932),
            .I(N__5925));
    InMux I__725 (
            .O(N__5931),
            .I(N__5922));
    LocalMux I__724 (
            .O(N__5928),
            .I(N__5917));
    Span4Mux_v I__723 (
            .O(N__5925),
            .I(N__5917));
    LocalMux I__722 (
            .O(N__5922),
            .I(\Lab_UT.secuu0.l_countZ0Z_5 ));
    Odrv4 I__721 (
            .O(N__5917),
            .I(\Lab_UT.secuu0.l_countZ0Z_5 ));
    CascadeMux I__720 (
            .O(N__5912),
            .I(N__5907));
    InMux I__719 (
            .O(N__5911),
            .I(N__5902));
    InMux I__718 (
            .O(N__5910),
            .I(N__5902));
    InMux I__717 (
            .O(N__5907),
            .I(N__5899));
    LocalMux I__716 (
            .O(N__5902),
            .I(\Lab_UT.secuu0.l_precountZ0Z_3 ));
    LocalMux I__715 (
            .O(N__5899),
            .I(\Lab_UT.secuu0.l_precountZ0Z_3 ));
    InMux I__714 (
            .O(N__5894),
            .I(N__5887));
    InMux I__713 (
            .O(N__5893),
            .I(N__5887));
    InMux I__712 (
            .O(N__5892),
            .I(N__5884));
    LocalMux I__711 (
            .O(N__5887),
            .I(\Lab_UT.secuu0.l_countZ0Z_15 ));
    LocalMux I__710 (
            .O(N__5884),
            .I(\Lab_UT.secuu0.l_countZ0Z_15 ));
    CascadeMux I__709 (
            .O(N__5879),
            .I(\Lab_UT.secuu0.un4_l_count_11_cascade_ ));
    InMux I__708 (
            .O(N__5876),
            .I(N__5863));
    InMux I__707 (
            .O(N__5875),
            .I(N__5863));
    InMux I__706 (
            .O(N__5874),
            .I(N__5863));
    InMux I__705 (
            .O(N__5873),
            .I(N__5863));
    InMux I__704 (
            .O(N__5872),
            .I(N__5860));
    LocalMux I__703 (
            .O(N__5863),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__702 (
            .O(N__5860),
            .I(\uu2.l_countZ0Z_1 ));
    CascadeMux I__701 (
            .O(N__5855),
            .I(N__5852));
    InMux I__700 (
            .O(N__5852),
            .I(N__5847));
    InMux I__699 (
            .O(N__5851),
            .I(N__5842));
    InMux I__698 (
            .O(N__5850),
            .I(N__5842));
    LocalMux I__697 (
            .O(N__5847),
            .I(N__5839));
    LocalMux I__696 (
            .O(N__5842),
            .I(\uu2.l_countZ0Z_3 ));
    Odrv12 I__695 (
            .O(N__5839),
            .I(\uu2.l_countZ0Z_3 ));
    CascadeMux I__694 (
            .O(N__5834),
            .I(\uu2.un3_r_clk_en_6_cascade_ ));
    CascadeMux I__693 (
            .O(N__5831),
            .I(uu2_un3_r_clk_en_0_cascade_));
    CEMux I__692 (
            .O(N__5828),
            .I(N__5824));
    SRMux I__691 (
            .O(N__5827),
            .I(N__5821));
    LocalMux I__690 (
            .O(N__5824),
            .I(N__5818));
    LocalMux I__689 (
            .O(N__5821),
            .I(N__5809));
    Span4Mux_s3_h I__688 (
            .O(N__5818),
            .I(N__5806));
    InMux I__687 (
            .O(N__5817),
            .I(N__5793));
    InMux I__686 (
            .O(N__5816),
            .I(N__5793));
    InMux I__685 (
            .O(N__5815),
            .I(N__5793));
    InMux I__684 (
            .O(N__5814),
            .I(N__5793));
    InMux I__683 (
            .O(N__5813),
            .I(N__5793));
    InMux I__682 (
            .O(N__5812),
            .I(N__5793));
    Span4Mux_s3_h I__681 (
            .O(N__5809),
            .I(N__5788));
    Span4Mux_h I__680 (
            .O(N__5806),
            .I(N__5788));
    LocalMux I__679 (
            .O(N__5793),
            .I(N__5785));
    Odrv4 I__678 (
            .O(N__5788),
            .I(\uu2.vbuf_tx_data_rdy ));
    Odrv4 I__677 (
            .O(N__5785),
            .I(\uu2.vbuf_tx_data_rdy ));
    InMux I__676 (
            .O(N__5780),
            .I(N__5777));
    LocalMux I__675 (
            .O(N__5777),
            .I(\uu2.un3_r_clk_en_0_0 ));
    CascadeMux I__674 (
            .O(N__5774),
            .I(N__5769));
    InMux I__673 (
            .O(N__5773),
            .I(N__5761));
    InMux I__672 (
            .O(N__5772),
            .I(N__5761));
    InMux I__671 (
            .O(N__5769),
            .I(N__5761));
    InMux I__670 (
            .O(N__5768),
            .I(N__5758));
    LocalMux I__669 (
            .O(N__5761),
            .I(\uu2.l_countZ0Z_2 ));
    LocalMux I__668 (
            .O(N__5758),
            .I(\uu2.l_countZ0Z_2 ));
    CascadeMux I__667 (
            .O(N__5753),
            .I(N__5749));
    CascadeMux I__666 (
            .O(N__5752),
            .I(N__5746));
    InMux I__665 (
            .O(N__5749),
            .I(N__5739));
    InMux I__664 (
            .O(N__5746),
            .I(N__5730));
    InMux I__663 (
            .O(N__5745),
            .I(N__5730));
    InMux I__662 (
            .O(N__5744),
            .I(N__5730));
    InMux I__661 (
            .O(N__5743),
            .I(N__5730));
    InMux I__660 (
            .O(N__5742),
            .I(N__5727));
    LocalMux I__659 (
            .O(N__5739),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__658 (
            .O(N__5730),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__657 (
            .O(N__5727),
            .I(\uu2.l_countZ0Z_0 ));
    InMux I__656 (
            .O(N__5720),
            .I(N__5717));
    LocalMux I__655 (
            .O(N__5717),
            .I(\uu2.un3_r_clk_en_7 ));
    InMux I__654 (
            .O(N__5714),
            .I(N__5711));
    LocalMux I__653 (
            .O(N__5711),
            .I(N__5708));
    Odrv4 I__652 (
            .O(N__5708),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__651 (
            .O(N__5705),
            .I(N__5702));
    LocalMux I__650 (
            .O(N__5702),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CascadeMux I__649 (
            .O(N__5699),
            .I(\uu2.un372_ci_cascade_ ));
    InMux I__648 (
            .O(N__5696),
            .I(N__5692));
    InMux I__647 (
            .O(N__5695),
            .I(N__5689));
    LocalMux I__646 (
            .O(N__5692),
            .I(\uu2.l_countZ0Z_10 ));
    LocalMux I__645 (
            .O(N__5689),
            .I(\uu2.l_countZ0Z_10 ));
    CascadeMux I__644 (
            .O(N__5684),
            .I(\uu2.un306_ci_cascade_ ));
    InMux I__643 (
            .O(N__5681),
            .I(N__5678));
    LocalMux I__642 (
            .O(N__5678),
            .I(\uu2.un339_ci_0 ));
    CascadeMux I__641 (
            .O(N__5675),
            .I(N__5672));
    InMux I__640 (
            .O(N__5672),
            .I(N__5668));
    CascadeMux I__639 (
            .O(N__5671),
            .I(N__5664));
    LocalMux I__638 (
            .O(N__5668),
            .I(N__5659));
    InMux I__637 (
            .O(N__5667),
            .I(N__5656));
    InMux I__636 (
            .O(N__5664),
            .I(N__5651));
    InMux I__635 (
            .O(N__5663),
            .I(N__5651));
    InMux I__634 (
            .O(N__5662),
            .I(N__5648));
    Odrv4 I__633 (
            .O(N__5659),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__632 (
            .O(N__5656),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__631 (
            .O(N__5651),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__630 (
            .O(N__5648),
            .I(\uu2.r_addrZ0Z_1 ));
    CascadeMux I__629 (
            .O(N__5639),
            .I(N__5636));
    InMux I__628 (
            .O(N__5636),
            .I(N__5633));
    LocalMux I__627 (
            .O(N__5633),
            .I(N__5627));
    InMux I__626 (
            .O(N__5632),
            .I(N__5624));
    InMux I__625 (
            .O(N__5631),
            .I(N__5621));
    InMux I__624 (
            .O(N__5630),
            .I(N__5618));
    Odrv4 I__623 (
            .O(N__5627),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__622 (
            .O(N__5624),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__621 (
            .O(N__5621),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__620 (
            .O(N__5618),
            .I(\uu2.r_addrZ0Z_2 ));
    CascadeMux I__619 (
            .O(N__5609),
            .I(N__5604));
    CascadeMux I__618 (
            .O(N__5608),
            .I(N__5601));
    CascadeMux I__617 (
            .O(N__5607),
            .I(N__5598));
    InMux I__616 (
            .O(N__5604),
            .I(N__5595));
    InMux I__615 (
            .O(N__5601),
            .I(N__5592));
    InMux I__614 (
            .O(N__5598),
            .I(N__5589));
    LocalMux I__613 (
            .O(N__5595),
            .I(N__5586));
    LocalMux I__612 (
            .O(N__5592),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__611 (
            .O(N__5589),
            .I(\uu2.r_addrZ0Z_3 ));
    Odrv4 I__610 (
            .O(N__5586),
            .I(\uu2.r_addrZ0Z_3 ));
    CascadeMux I__609 (
            .O(N__5579),
            .I(N__5576));
    InMux I__608 (
            .O(N__5576),
            .I(N__5573));
    LocalMux I__607 (
            .O(N__5573),
            .I(N__5569));
    InMux I__606 (
            .O(N__5572),
            .I(N__5562));
    Span12Mux_s3_h I__605 (
            .O(N__5569),
            .I(N__5559));
    InMux I__604 (
            .O(N__5568),
            .I(N__5556));
    InMux I__603 (
            .O(N__5567),
            .I(N__5549));
    InMux I__602 (
            .O(N__5566),
            .I(N__5549));
    InMux I__601 (
            .O(N__5565),
            .I(N__5549));
    LocalMux I__600 (
            .O(N__5562),
            .I(N__5546));
    Odrv12 I__599 (
            .O(N__5559),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__598 (
            .O(N__5556),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__597 (
            .O(N__5549),
            .I(\uu2.r_addrZ0Z_0 ));
    Odrv4 I__596 (
            .O(N__5546),
            .I(\uu2.r_addrZ0Z_0 ));
    InMux I__595 (
            .O(N__5537),
            .I(N__5526));
    InMux I__594 (
            .O(N__5536),
            .I(N__5526));
    InMux I__593 (
            .O(N__5535),
            .I(N__5526));
    InMux I__592 (
            .O(N__5534),
            .I(N__5521));
    InMux I__591 (
            .O(N__5533),
            .I(N__5521));
    LocalMux I__590 (
            .O(N__5526),
            .I(N__5518));
    LocalMux I__589 (
            .O(N__5521),
            .I(\uu2.un415_ci_0 ));
    Odrv4 I__588 (
            .O(N__5518),
            .I(\uu2.un415_ci_0 ));
    CascadeMux I__587 (
            .O(N__5513),
            .I(\uu2.vbuf_raddr.un459_ci_0_cascade_ ));
    CascadeMux I__586 (
            .O(N__5510),
            .I(N__5507));
    InMux I__585 (
            .O(N__5507),
            .I(N__5503));
    InMux I__584 (
            .O(N__5506),
            .I(N__5500));
    LocalMux I__583 (
            .O(N__5503),
            .I(\uu2.r_addrZ0Z_8 ));
    LocalMux I__582 (
            .O(N__5500),
            .I(\uu2.r_addrZ0Z_8 ));
    CascadeMux I__581 (
            .O(N__5495),
            .I(N__5491));
    CascadeMux I__580 (
            .O(N__5494),
            .I(N__5488));
    InMux I__579 (
            .O(N__5491),
            .I(N__5483));
    InMux I__578 (
            .O(N__5488),
            .I(N__5476));
    InMux I__577 (
            .O(N__5487),
            .I(N__5476));
    InMux I__576 (
            .O(N__5486),
            .I(N__5476));
    LocalMux I__575 (
            .O(N__5483),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__574 (
            .O(N__5476),
            .I(\uu2.r_addrZ0Z_6 ));
    CascadeMux I__573 (
            .O(N__5471),
            .I(N__5468));
    InMux I__572 (
            .O(N__5468),
            .I(N__5463));
    InMux I__571 (
            .O(N__5467),
            .I(N__5458));
    InMux I__570 (
            .O(N__5466),
            .I(N__5458));
    LocalMux I__569 (
            .O(N__5463),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__568 (
            .O(N__5458),
            .I(\uu2.r_addrZ0Z_7 ));
    CascadeMux I__567 (
            .O(N__5453),
            .I(N__5450));
    InMux I__566 (
            .O(N__5450),
            .I(N__5447));
    LocalMux I__565 (
            .O(N__5447),
            .I(N__5441));
    InMux I__564 (
            .O(N__5446),
            .I(N__5438));
    InMux I__563 (
            .O(N__5445),
            .I(N__5435));
    InMux I__562 (
            .O(N__5444),
            .I(N__5432));
    Odrv4 I__561 (
            .O(N__5441),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__560 (
            .O(N__5438),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__559 (
            .O(N__5435),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__558 (
            .O(N__5432),
            .I(\uu2.r_addrZ0Z_5 ));
    CascadeMux I__557 (
            .O(N__5423),
            .I(N__5420));
    InMux I__556 (
            .O(N__5420),
            .I(N__5416));
    CascadeMux I__555 (
            .O(N__5419),
            .I(N__5412));
    LocalMux I__554 (
            .O(N__5416),
            .I(N__5407));
    InMux I__553 (
            .O(N__5415),
            .I(N__5404));
    InMux I__552 (
            .O(N__5412),
            .I(N__5397));
    InMux I__551 (
            .O(N__5411),
            .I(N__5397));
    InMux I__550 (
            .O(N__5410),
            .I(N__5397));
    Odrv4 I__549 (
            .O(N__5407),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__548 (
            .O(N__5404),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__547 (
            .O(N__5397),
            .I(\uu2.r_addrZ0Z_4 ));
    CascadeMux I__546 (
            .O(N__5390),
            .I(N__5387));
    InMux I__545 (
            .O(N__5387),
            .I(N__5381));
    InMux I__544 (
            .O(N__5386),
            .I(N__5381));
    LocalMux I__543 (
            .O(N__5381),
            .I(\uu2.vbuf_raddr.un437_ci_3 ));
    CascadeMux I__542 (
            .O(N__5378),
            .I(\uu2.mem0.g0_0_a3_3_cascade_ ));
    InMux I__541 (
            .O(N__5375),
            .I(N__5372));
    LocalMux I__540 (
            .O(N__5372),
            .I(\uu2.mem0.w_data_1 ));
    CascadeMux I__539 (
            .O(N__5369),
            .I(\uu2.mem0.g1_0_6_cascade_ ));
    InMux I__538 (
            .O(N__5366),
            .I(N__5363));
    LocalMux I__537 (
            .O(N__5363),
            .I(\uu2.mem0.N_4_i ));
    CascadeMux I__536 (
            .O(N__5360),
            .I(N__5357));
    InMux I__535 (
            .O(N__5357),
            .I(N__5354));
    LocalMux I__534 (
            .O(N__5354),
            .I(\uu2.mem0.w_addr_6 ));
    InMux I__533 (
            .O(N__5351),
            .I(N__5348));
    LocalMux I__532 (
            .O(N__5348),
            .I(\uu2.mem0.N_14_0 ));
    InMux I__531 (
            .O(N__5345),
            .I(N__5342));
    LocalMux I__530 (
            .O(N__5342),
            .I(\Lab_UT.secuu0.un208_ci_0 ));
    InMux I__529 (
            .O(N__5339),
            .I(N__5333));
    InMux I__528 (
            .O(N__5338),
            .I(N__5333));
    LocalMux I__527 (
            .O(N__5333),
            .I(\Lab_UT.secuu0.l_countZ0Z_13 ));
    InMux I__526 (
            .O(N__5330),
            .I(N__5324));
    InMux I__525 (
            .O(N__5329),
            .I(N__5321));
    InMux I__524 (
            .O(N__5328),
            .I(N__5318));
    InMux I__523 (
            .O(N__5327),
            .I(N__5315));
    LocalMux I__522 (
            .O(N__5324),
            .I(\Lab_UT.secuu0.l_countZ0Z_10 ));
    LocalMux I__521 (
            .O(N__5321),
            .I(\Lab_UT.secuu0.l_countZ0Z_10 ));
    LocalMux I__520 (
            .O(N__5318),
            .I(\Lab_UT.secuu0.l_countZ0Z_10 ));
    LocalMux I__519 (
            .O(N__5315),
            .I(\Lab_UT.secuu0.l_countZ0Z_10 ));
    InMux I__518 (
            .O(N__5306),
            .I(N__5294));
    InMux I__517 (
            .O(N__5305),
            .I(N__5294));
    InMux I__516 (
            .O(N__5304),
            .I(N__5294));
    InMux I__515 (
            .O(N__5303),
            .I(N__5287));
    InMux I__514 (
            .O(N__5302),
            .I(N__5287));
    InMux I__513 (
            .O(N__5301),
            .I(N__5287));
    LocalMux I__512 (
            .O(N__5294),
            .I(\Lab_UT.secuu0.l_countZ0Z_8 ));
    LocalMux I__511 (
            .O(N__5287),
            .I(\Lab_UT.secuu0.l_countZ0Z_8 ));
    CascadeMux I__510 (
            .O(N__5282),
            .I(N__5279));
    InMux I__509 (
            .O(N__5279),
            .I(N__5276));
    LocalMux I__508 (
            .O(N__5276),
            .I(\uu2.mem0.w_addr_8 ));
    CascadeMux I__507 (
            .O(N__5273),
            .I(N__5270));
    InMux I__506 (
            .O(N__5270),
            .I(N__5267));
    LocalMux I__505 (
            .O(N__5267),
            .I(\uu2.mem0.w_addr_1 ));
    CascadeMux I__504 (
            .O(N__5264),
            .I(N__5261));
    InMux I__503 (
            .O(N__5261),
            .I(N__5258));
    LocalMux I__502 (
            .O(N__5258),
            .I(N__5255));
    Odrv4 I__501 (
            .O(N__5255),
            .I(\uu2.mem0.w_addr_2 ));
    CascadeMux I__500 (
            .O(N__5252),
            .I(N__5249));
    InMux I__499 (
            .O(N__5249),
            .I(N__5246));
    LocalMux I__498 (
            .O(N__5246),
            .I(\uu2.mem0.w_addr_5 ));
    InMux I__497 (
            .O(N__5243),
            .I(N__5240));
    LocalMux I__496 (
            .O(N__5240),
            .I(\uu2.mem0.w_data_4 ));
    CascadeMux I__495 (
            .O(N__5237),
            .I(N__5234));
    InMux I__494 (
            .O(N__5234),
            .I(N__5231));
    LocalMux I__493 (
            .O(N__5231),
            .I(\uu2.mem0.w_addr_3 ));
    CascadeMux I__492 (
            .O(N__5228),
            .I(\Lab_UT.secuu0.un230_ci_1_cascade_ ));
    CascadeMux I__491 (
            .O(N__5225),
            .I(N__5219));
    CascadeMux I__490 (
            .O(N__5224),
            .I(N__5216));
    CascadeMux I__489 (
            .O(N__5223),
            .I(N__5211));
    InMux I__488 (
            .O(N__5222),
            .I(N__5208));
    InMux I__487 (
            .O(N__5219),
            .I(N__5197));
    InMux I__486 (
            .O(N__5216),
            .I(N__5197));
    InMux I__485 (
            .O(N__5215),
            .I(N__5197));
    InMux I__484 (
            .O(N__5214),
            .I(N__5197));
    InMux I__483 (
            .O(N__5211),
            .I(N__5197));
    LocalMux I__482 (
            .O(N__5208),
            .I(N__5194));
    LocalMux I__481 (
            .O(N__5197),
            .I(\Lab_UT.secuu0.l_precountZ0Z_0 ));
    Odrv4 I__480 (
            .O(N__5194),
            .I(\Lab_UT.secuu0.l_precountZ0Z_0 ));
    InMux I__479 (
            .O(N__5189),
            .I(N__5185));
    InMux I__478 (
            .O(N__5188),
            .I(N__5182));
    LocalMux I__477 (
            .O(N__5185),
            .I(N__5178));
    LocalMux I__476 (
            .O(N__5182),
            .I(N__5174));
    InMux I__475 (
            .O(N__5181),
            .I(N__5171));
    Span4Mux_s3_h I__474 (
            .O(N__5178),
            .I(N__5168));
    InMux I__473 (
            .O(N__5177),
            .I(N__5165));
    Odrv4 I__472 (
            .O(N__5174),
            .I(\Lab_UT.secuu0.l_countZ0Z_4 ));
    LocalMux I__471 (
            .O(N__5171),
            .I(\Lab_UT.secuu0.l_countZ0Z_4 ));
    Odrv4 I__470 (
            .O(N__5168),
            .I(\Lab_UT.secuu0.l_countZ0Z_4 ));
    LocalMux I__469 (
            .O(N__5165),
            .I(\Lab_UT.secuu0.l_countZ0Z_4 ));
    CascadeMux I__468 (
            .O(N__5156),
            .I(\Lab_UT.secuu0.un4_l_count_14_cascade_ ));
    InMux I__467 (
            .O(N__5153),
            .I(N__5146));
    InMux I__466 (
            .O(N__5152),
            .I(N__5146));
    InMux I__465 (
            .O(N__5151),
            .I(N__5143));
    LocalMux I__464 (
            .O(N__5146),
            .I(\Lab_UT.secuu0.un4_l_count_0_8 ));
    LocalMux I__463 (
            .O(N__5143),
            .I(\Lab_UT.secuu0.un4_l_count_0_8 ));
    CascadeMux I__462 (
            .O(N__5138),
            .I(\Lab_UT.secuu0.un4_l_count_0_8_cascade_ ));
    CascadeMux I__461 (
            .O(N__5135),
            .I(N__5129));
    InMux I__460 (
            .O(N__5134),
            .I(N__5124));
    InMux I__459 (
            .O(N__5133),
            .I(N__5124));
    InMux I__458 (
            .O(N__5132),
            .I(N__5119));
    InMux I__457 (
            .O(N__5129),
            .I(N__5119));
    LocalMux I__456 (
            .O(N__5124),
            .I(\Lab_UT.secuu0.l_countZ0Z_14 ));
    LocalMux I__455 (
            .O(N__5119),
            .I(\Lab_UT.secuu0.l_countZ0Z_14 ));
    InMux I__454 (
            .O(N__5114),
            .I(N__5106));
    InMux I__453 (
            .O(N__5113),
            .I(N__5106));
    InMux I__452 (
            .O(N__5112),
            .I(N__5101));
    InMux I__451 (
            .O(N__5111),
            .I(N__5101));
    LocalMux I__450 (
            .O(N__5106),
            .I(\Lab_UT.secuu0.un197_ci_9 ));
    LocalMux I__449 (
            .O(N__5101),
            .I(\Lab_UT.secuu0.un197_ci_9 ));
    CascadeMux I__448 (
            .O(N__5096),
            .I(N__5093));
    InMux I__447 (
            .O(N__5093),
            .I(N__5088));
    InMux I__446 (
            .O(N__5092),
            .I(N__5085));
    InMux I__445 (
            .O(N__5091),
            .I(N__5082));
    LocalMux I__444 (
            .O(N__5088),
            .I(\Lab_UT.secuu0.l_countZ0Z_12 ));
    LocalMux I__443 (
            .O(N__5085),
            .I(\Lab_UT.secuu0.l_countZ0Z_12 ));
    LocalMux I__442 (
            .O(N__5082),
            .I(\Lab_UT.secuu0.l_countZ0Z_12 ));
    CascadeMux I__441 (
            .O(N__5075),
            .I(\Lab_UT.secuu0.un197_ci_9_cascade_ ));
    IoInMux I__440 (
            .O(N__5072),
            .I(N__5069));
    LocalMux I__439 (
            .O(N__5069),
            .I(\resetGen.rst_isoZ0 ));
    CascadeMux I__438 (
            .O(N__5066),
            .I(\Lab_UT.secuu0.un131_ci_3_cascade_ ));
    InMux I__437 (
            .O(N__5063),
            .I(N__5060));
    LocalMux I__436 (
            .O(N__5060),
            .I(N__5057));
    Odrv4 I__435 (
            .O(N__5057),
            .I(uart_RXD));
    IoInMux I__434 (
            .O(N__5054),
            .I(N__5051));
    LocalMux I__433 (
            .O(N__5051),
            .I(N__5048));
    IoSpan4Mux I__432 (
            .O(N__5048),
            .I(N__5045));
    Odrv4 I__431 (
            .O(N__5045),
            .I(clk_in_c));
    INV \INVuu2.w_addr_displaying_fast_5C  (
            .O(\INVuu2.w_addr_displaying_fast_5C_net ),
            .I(N__13408));
    INV \INVuu2.w_addr_displaying_8C  (
            .O(\INVuu2.w_addr_displaying_8C_net ),
            .I(N__13396));
    INV \INVuu2.w_addr_displaying_fast_1C  (
            .O(\INVuu2.w_addr_displaying_fast_1C_net ),
            .I(N__13401));
    INV \INVuu2.w_addr_displaying_fast_0C  (
            .O(\INVuu2.w_addr_displaying_fast_0C_net ),
            .I(N__13407));
    INV \INVuu2.w_addr_displaying_fast_6C  (
            .O(\INVuu2.w_addr_displaying_fast_6C_net ),
            .I(N__13413));
    INV \INVuu2.w_addr_user_0C  (
            .O(\INVuu2.w_addr_user_0C_net ),
            .I(N__13430));
    INV \INVuu2.w_addr_displaying_3_rep1C  (
            .O(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .I(N__13390));
    INV \INVuu2.w_addr_displaying_0_rep1C  (
            .O(\INVuu2.w_addr_displaying_0_rep1C_net ),
            .I(N__13395));
    INV \INVuu2.w_addr_displaying_2_rep1C  (
            .O(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .I(N__13400));
    INV \INVuu2.w_addr_displaying_5_rep1C  (
            .O(\INVuu2.w_addr_displaying_5_rep1C_net ),
            .I(N__13406));
    INV \INVuu2.w_addr_user_5C  (
            .O(\INVuu2.w_addr_user_5C_net ),
            .I(N__13412));
    INV \INVuu2.w_addr_user_7C  (
            .O(\INVuu2.w_addr_user_7C_net ),
            .I(N__13417));
    INV \INVuu2.w_addr_user_2C  (
            .O(\INVuu2.w_addr_user_2C_net ),
            .I(N__13424));
    INV \INVuu2.w_addr_displaying_8_rep1C  (
            .O(\INVuu2.w_addr_displaying_8_rep1C_net ),
            .I(N__13383));
    INV \INVuu2.w_addr_displaying_5C  (
            .O(\INVuu2.w_addr_displaying_5C_net ),
            .I(N__13397));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_12_0_));
    ICE_GB \resetGen.rst_iso_RNIEOGF  (
            .USERSIGNALTOGLOBALBUFFER(N__5072),
            .GLOBALBUFFEROUTPUT(resetGen_rst_iso_g));
    ICE_GB \Lab_UT.secuu0.delay_line_RNILBAI7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__6314),
            .GLOBALBUFFEROUTPUT(\Lab_UT.secuu0.un11_l_count_i_g ));
    ICE_GB \latticehx1k_pll_inst.PLLOUTCORE_derived_clock_RNIALC1  (
            .USERSIGNALTOGLOBALBUFFER(N__7613),
            .GLOBALBUFFEROUTPUT(clk_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \resetGen.rst_iso_LC_1_8_0 .C_ON=1'b0;
    defparam \resetGen.rst_iso_LC_1_8_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_iso_LC_1_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_iso_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6728),
            .lcout(\resetGen.rst_isoZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13426),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_5_LC_2_5_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_5_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_5_LC_2_5_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \Lab_UT.secuu0.l_count_5_LC_2_5_0  (
            .in0(N__6425),
            .in1(N__5188),
            .in2(_gnd_net_),
            .in3(N__5935),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13432),
            .ce(N__6370),
            .sr(N__12307));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_3_LC_2_6_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_3_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_3_LC_2_6_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_3_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__5931),
            .in2(_gnd_net_),
            .in3(N__5189),
            .lcout(\Lab_UT.secuu0.un131_ci_3 ),
            .ltout(\Lab_UT.secuu0.un131_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_7__un142_ci_0_LC_2_6_2 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_7__un142_ci_0_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_7__un142_ci_0_LC_2_6_2 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_7__un142_ci_0_LC_2_6_2  (
            .in0(_gnd_net_),
            .in1(N__6518),
            .in2(N__5066),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.secuu0.un142_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_0_LC_2_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.hh_0_LC_2_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_2_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5063),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13404),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.sec_clk_LC_4_4_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.sec_clk_LC_4_4_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.sec_clk_LC_4_4_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.secuu0.sec_clk_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__6464),
            .in2(_gnd_net_),
            .in3(N__13107),
            .lcout(Lab_UT_l_oneSecPluse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13429),
            .ce(),
            .sr(N__12311));
    defparam \Lab_UT.secuu0.delay_line_1_LC_4_4_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.delay_line_1_LC_4_4_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.delay_line_1_LC_4_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.secuu0.delay_line_1_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6326),
            .lcout(\Lab_UT.secuu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13429),
            .ce(),
            .sr(N__12311));
    defparam \Lab_UT.secuu0.l_precount_0_LC_4_4_2 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_precount_0_LC_4_4_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_precount_0_LC_4_4_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.secuu0.l_precount_0_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5214),
            .lcout(\Lab_UT.secuu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13429),
            .ce(),
            .sr(N__12311));
    defparam \Lab_UT.secuu0.l_precount_3_LC_4_4_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_precount_3_LC_4_4_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_precount_3_LC_4_4_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \Lab_UT.secuu0.l_precount_3_LC_4_4_3  (
            .in0(N__5977),
            .in1(N__5911),
            .in2(N__5225),
            .in3(N__5957),
            .lcout(\Lab_UT.secuu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13429),
            .ce(),
            .sr(N__12311));
    defparam \Lab_UT.secuu0.l_precount_2_LC_4_4_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_precount_2_LC_4_4_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_precount_2_LC_4_4_5 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \Lab_UT.secuu0.l_precount_2_LC_4_4_5  (
            .in0(N__5976),
            .in1(_gnd_net_),
            .in2(N__5224),
            .in3(N__5956),
            .lcout(\Lab_UT.secuu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13429),
            .ce(),
            .sr(N__12311));
    defparam \Lab_UT.secuu0.l_precount_1_LC_4_4_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_precount_1_LC_4_4_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_precount_1_LC_4_4_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.secuu0.l_precount_1_LC_4_4_6  (
            .in0(N__5955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5215),
            .lcout(\Lab_UT.secuu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13429),
            .ce(),
            .sr(N__12311));
    defparam \Lab_UT.secuu0.delay_line_0_LC_4_4_7 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.delay_line_0_LC_4_4_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.delay_line_0_LC_4_4_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.delay_line_0_LC_4_4_7  (
            .in0(N__5975),
            .in1(N__5910),
            .in2(N__5223),
            .in3(N__5954),
            .lcout(\Lab_UT.secuu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13429),
            .ce(),
            .sr(N__12311));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_13__un208_ci_0_LC_4_5_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_13__un208_ci_0_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_13__un208_ci_0_LC_4_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_13__un208_ci_0_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(N__5111),
            .in2(_gnd_net_),
            .in3(N__5092),
            .lcout(\Lab_UT.secuu0.un208_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_11__un186_ci_0_LC_4_5_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_11__un186_ci_0_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_11__un186_ci_0_LC_4_5_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_11__un186_ci_0_LC_4_5_1  (
            .in0(N__5305),
            .in1(N__6212),
            .in2(_gnd_net_),
            .in3(N__5329),
            .lcout(\Lab_UT.secuu0.un186_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_12__un197_ci_9_LC_4_5_2 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_12__un197_ci_9_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_12__un197_ci_9_LC_4_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_12__un197_ci_9_LC_4_5_2  (
            .in0(N__6286),
            .in1(N__5328),
            .in2(N__6217),
            .in3(N__5304),
            .lcout(\Lab_UT.secuu0.un197_ci_9 ),
            .ltout(\Lab_UT.secuu0.un197_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_16__un241_ci_2_LC_4_5_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_16__un241_ci_2_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_16__un241_ci_2_LC_4_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_16__un241_ci_2_LC_4_5_3  (
            .in0(N__5893),
            .in1(N__5133),
            .in2(N__5075),
            .in3(N__5152),
            .lcout(\Lab_UT.secuu0.un241_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_9_LC_4_5_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_9_LC_4_5_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_9_LC_4_5_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \Lab_UT.secuu0.l_count_9_LC_4_5_4  (
            .in0(N__6213),
            .in1(N__6582),
            .in2(_gnd_net_),
            .in3(N__5306),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13427),
            .ce(N__6372),
            .sr(N__12309));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_15__un230_ci_1_LC_4_5_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_15__un230_ci_1_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_15__un230_ci_1_LC_4_5_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_15__un230_ci_1_LC_4_5_5  (
            .in0(N__5112),
            .in1(N__5134),
            .in2(_gnd_net_),
            .in3(N__5153),
            .lcout(),
            .ltout(\Lab_UT.secuu0.un230_ci_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_15_LC_4_5_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_15_LC_4_5_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_15_LC_4_5_6 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \Lab_UT.secuu0.l_count_15_LC_4_5_6  (
            .in0(N__6581),
            .in1(N__6485),
            .in2(N__5228),
            .in3(N__5894),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13427),
            .ce(N__6372),
            .sr(N__12309));
    defparam \Lab_UT.secuu0.l_count_4_LC_4_5_7 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_4_LC_4_5_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_4_LC_4_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Lab_UT.secuu0.l_count_4_LC_4_5_7  (
            .in0(N__6486),
            .in1(N__6417),
            .in2(_gnd_net_),
            .in3(N__5181),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13427),
            .ce(N__6372),
            .sr(N__12309));
    defparam \Lab_UT.secuu0.l_count_RNI0S951_2_LC_4_6_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNI0S951_2_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNI0S951_2_LC_4_6_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.secuu0.l_count_RNI0S951_2_LC_4_6_0  (
            .in0(N__5327),
            .in1(N__5301),
            .in2(N__5135),
            .in3(N__6650),
            .lcout(),
            .ltout(\Lab_UT.secuu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_RNI20OC2_4_LC_4_6_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNI20OC2_4_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNI20OC2_4_LC_4_6_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNI20OC2_4_LC_4_6_1  (
            .in0(N__5222),
            .in1(N__5177),
            .in2(N__5156),
            .in3(N__5151),
            .lcout(\Lab_UT.secuu0.un4_l_count_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_RNIFM2M_13_LC_4_6_2 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNIFM2M_13_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNIFM2M_13_LC_4_6_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNIFM2M_13_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__5338),
            .in2(_gnd_net_),
            .in3(N__5091),
            .lcout(\Lab_UT.secuu0.un4_l_count_0_8 ),
            .ltout(\Lab_UT.secuu0.un4_l_count_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_14_LC_4_6_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_14_LC_4_6_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_14_LC_4_6_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \Lab_UT.secuu0.l_count_14_LC_4_6_3  (
            .in0(N__5114),
            .in1(N__6575),
            .in2(N__5138),
            .in3(N__5132),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13422),
            .ce(N__6371),
            .sr(N__12308));
    defparam \Lab_UT.secuu0.l_count_12_LC_4_6_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_12_LC_4_6_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_12_LC_4_6_4 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \Lab_UT.secuu0.l_count_12_LC_4_6_4  (
            .in0(N__6573),
            .in1(N__6487),
            .in2(N__5096),
            .in3(N__5113),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13422),
            .ce(N__6371),
            .sr(N__12308));
    defparam \Lab_UT.secuu0.l_count_13_LC_4_6_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_13_LC_4_6_5 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_13_LC_4_6_5 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \Lab_UT.secuu0.l_count_13_LC_4_6_5  (
            .in0(N__5339),
            .in1(N__5345),
            .in2(N__6491),
            .in3(N__6574),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13422),
            .ce(N__6371),
            .sr(N__12308));
    defparam \Lab_UT.secuu0.l_count_10_LC_4_6_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_10_LC_4_6_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_10_LC_4_6_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \Lab_UT.secuu0.l_count_10_LC_4_6_6  (
            .in0(N__6576),
            .in1(N__5330),
            .in2(N__6218),
            .in3(N__5302),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13422),
            .ce(N__6371),
            .sr(N__12308));
    defparam \Lab_UT.secuu0.l_count_8_LC_4_6_7 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_8_LC_4_6_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_8_LC_4_6_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.secuu0.l_count_8_LC_4_6_7  (
            .in0(N__5303),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6572),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13422),
            .ce(N__6371),
            .sr(N__12308));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_7_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_4_7_1  (
            .in0(N__11248),
            .in1(N__8171),
            .in2(_gnd_net_),
            .in3(N__9967),
            .lcout(\uu2.mem0.w_addr_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_7_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_4_7_2  (
            .in0(N__7934),
            .in1(N__11249),
            .in2(_gnd_net_),
            .in3(N__11694),
            .lcout(\uu2.mem0.w_addr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_4_7_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_4_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_4_7_3  (
            .in0(N__11245),
            .in1(N__8120),
            .in2(_gnd_net_),
            .in3(N__11596),
            .lcout(\uu2.mem0.w_addr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_4_7_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_4_7_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_4_7_5  (
            .in0(N__11247),
            .in1(_gnd_net_),
            .in2(N__8033),
            .in3(N__11872),
            .lcout(\uu2.mem0.w_addr_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_7_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_7_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_4_7_6  (
            .in0(N__10967),
            .in1(N__6857),
            .in2(_gnd_net_),
            .in3(N__11250),
            .lcout(\uu2.mem0.w_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_7_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_4_7_7  (
            .in0(N__11246),
            .in1(N__7808),
            .in2(_gnd_net_),
            .in3(N__12079),
            .lcout(\uu2.mem0.w_addr_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_4_8_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_4_8_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_23_LC_4_8_0  (
            .in0(N__6890),
            .in1(N__5351),
            .in2(N__7022),
            .in3(N__6905),
            .lcout(),
            .ltout(\uu2.mem0.g0_0_a3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_8_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_8_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_4_8_1  (
            .in0(N__6821),
            .in1(N__6866),
            .in2(N__5378),
            .in3(N__5366),
            .lcout(\uu2.mem0.w_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_4_8_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_4_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_31_LC_4_8_2  (
            .in0(_gnd_net_),
            .in1(N__6884),
            .in2(_gnd_net_),
            .in3(N__6851),
            .lcout(),
            .ltout(\uu2.mem0.g1_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_4_8_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_4_8_3 .LUT_INIT=16'b0111010001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_19_LC_4_8_3  (
            .in0(N__6839),
            .in1(N__11251),
            .in2(N__5369),
            .in3(N__9707),
            .lcout(\uu2.mem0.N_4_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_4_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_4_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_4_8_4  (
            .in0(N__11252),
            .in1(N__8087),
            .in2(_gnd_net_),
            .in3(N__9865),
            .lcout(\uu2.mem0.w_addr_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_4_8_6 .C_ON=1'b0;
    defparam \resetGen.rst_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_4_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6713),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13410),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_4_8_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_4_8_7 .LUT_INIT=16'b0000110010001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_36_LC_4_8_7  (
            .in0(N__12077),
            .in1(N__8333),
            .in2(N__11597),
            .in3(N__8549),
            .lcout(\uu2.mem0.N_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_3_LC_4_9_0 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_4_9_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_4_9_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_4_9_0  (
            .in0(N__5632),
            .in1(N__5667),
            .in2(N__5607),
            .in3(N__5568),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13405),
            .ce(N__7246),
            .sr(N__12298));
    defparam \uu2.r_addr_esr_6_LC_4_9_1 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_4_9_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_4_9_1 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_6_LC_4_9_1  (
            .in0(N__5446),
            .in1(N__5415),
            .in2(N__5494),
            .in3(N__5535),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13405),
            .ce(N__7246),
            .sr(N__12298));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un459_ci_0_LC_4_9_2 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un459_ci_0_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un459_ci_0_LC_4_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un459_ci_0_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(N__5466),
            .in2(_gnd_net_),
            .in3(N__5486),
            .lcout(),
            .ltout(\uu2.vbuf_raddr.un459_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_8_LC_4_9_3 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_4_9_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_4_9_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_8_LC_4_9_3  (
            .in0(N__5506),
            .in1(N__5386),
            .in2(N__5513),
            .in3(N__5536),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13405),
            .ce(N__7246),
            .sr(N__12298));
    defparam \uu2.r_addr_esr_7_LC_4_9_4 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_4_9_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_4_9_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_7_LC_4_9_4  (
            .in0(N__5537),
            .in1(N__5467),
            .in2(N__5390),
            .in3(N__5487),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13405),
            .ce(N__7246),
            .sr(N__12298));
    defparam \uu2.r_addr_2_LC_4_10_0 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_4_10_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_4_10_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_2_LC_4_10_0  (
            .in0(N__5815),
            .in1(N__5631),
            .in2(N__5671),
            .in3(N__5567),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13398),
            .ce(),
            .sr(N__12322));
    defparam \uu2.r_addr_1_LC_4_10_1 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_4_10_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_4_10_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.r_addr_1_LC_4_10_1  (
            .in0(N__5566),
            .in1(N__5663),
            .in2(_gnd_net_),
            .in3(N__5816),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13398),
            .ce(),
            .sr(N__12322));
    defparam \uu2.r_addr_0_LC_4_10_2 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_4_10_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_4_10_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.r_addr_0_LC_4_10_2  (
            .in0(N__5813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5565),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13398),
            .ce(),
            .sr(N__12322));
    defparam \uu2.l_count_RNI88MU5_4_LC_4_10_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNI88MU5_4_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI88MU5_4_LC_4_10_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.l_count_RNI88MU5_4_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__12321),
            .in2(_gnd_net_),
            .in3(N__5812),
            .lcout(\uu2.vbuf_tx_data_rdy_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_4_LC_4_10_4 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_4_10_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_4_10_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.r_addr_4_LC_4_10_4  (
            .in0(N__5814),
            .in1(N__5411),
            .in2(_gnd_net_),
            .in3(N__5533),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13398),
            .ce(),
            .sr(N__12322));
    defparam \uu2.r_addr_5_LC_4_10_5 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_4_10_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_4_10_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_5_LC_4_10_5  (
            .in0(N__5534),
            .in1(N__5445),
            .in2(N__5419),
            .in3(N__5817),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13398),
            .ce(),
            .sr(N__12322));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un437_ci_3_LC_4_10_6 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un437_ci_3_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un437_ci_3_LC_4_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un437_ci_3_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(N__5444),
            .in2(_gnd_net_),
            .in3(N__5410),
            .lcout(\uu2.vbuf_raddr.un437_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_1_LC_4_11_0 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_4_11_0 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_1_LC_4_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_1_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(N__5745),
            .in2(_gnd_net_),
            .in3(N__5874),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13393),
            .ce(),
            .sr(N__12299));
    defparam \uu2.l_count_3_LC_4_11_1 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_4_11_1 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_3_LC_4_11_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.l_count_3_LC_4_11_1  (
            .in0(N__5876),
            .in1(N__5773),
            .in2(N__5752),
            .in3(N__5851),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13393),
            .ce(),
            .sr(N__12299));
    defparam \uu2.l_count_2_LC_4_11_2 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_2_LC_4_11_2 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \uu2.l_count_2_LC_4_11_2  (
            .in0(N__5772),
            .in1(N__10476),
            .in2(N__5753),
            .in3(N__5875),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13393),
            .ce(),
            .sr(N__12299));
    defparam \uu2.l_count_0_LC_4_11_3 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_4_11_3 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_0_LC_4_11_3 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \uu2.l_count_0_LC_4_11_3  (
            .in0(N__5744),
            .in1(_gnd_net_),
            .in2(N__10506),
            .in3(_gnd_net_),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13393),
            .ce(),
            .sr(N__12299));
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_11_4 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_11_4  (
            .in0(N__5850),
            .in1(N__5743),
            .in2(N__5774),
            .in3(N__5873),
            .lcout(\uu2.un306_ci ),
            .ltout(\uu2.un306_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_7_LC_4_11_5 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_7_LC_4_11_5 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu2.l_count_7_LC_4_11_5  (
            .in0(N__10472),
            .in1(N__5681),
            .in2(N__5684),
            .in3(N__6172),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13393),
            .ce(),
            .sr(N__12299));
    defparam \uu2.vbuf_count.counter_gen_label_7__un339_ci_0_LC_4_11_6 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_7__un339_ci_0_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_7__un339_ci_0_LC_4_11_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_7__un339_ci_0_LC_4_11_6  (
            .in0(N__6014),
            .in1(N__6098),
            .in2(_gnd_net_),
            .in3(N__6071),
            .lcout(\uu2.un339_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un415_ci_LC_4_11_7 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un415_ci_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un415_ci_LC_4_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un415_ci_LC_4_11_7  (
            .in0(N__5662),
            .in1(N__5630),
            .in2(N__5609),
            .in3(N__5572),
            .lcout(\uu2.un415_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_6_LC_4_12_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_6_LC_4_12_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \buart.Z_tx.shifter_6_LC_4_12_0  (
            .in0(N__10286),
            .in1(N__5714),
            .in2(N__10507),
            .in3(N__7058),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13388),
            .ce(N__8588),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNICDGK1_3_LC_4_12_1 .C_ON=1'b0;
    defparam \uu2.l_count_RNICDGK1_3_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNICDGK1_3_LC_4_12_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uu2.l_count_RNICDGK1_3_LC_4_12_1  (
            .in0(N__6168),
            .in1(N__5872),
            .in2(N__5855),
            .in3(N__6111),
            .lcout(),
            .ltout(\uu2.un3_r_clk_en_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI0NA44_4_LC_4_12_2 .C_ON=1'b0;
    defparam \uu2.l_count_RNI0NA44_4_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI0NA44_4_LC_4_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI0NA44_4_LC_4_12_2  (
            .in0(N__6013),
            .in1(N__5720),
            .in2(N__5834),
            .in3(N__5780),
            .lcout(uu2_un3_r_clk_en_0),
            .ltout(uu2_un3_r_clk_en_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIQF5F5_4_LC_4_12_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNIQF5F5_4_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIQF5F5_4_LC_4_12_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.l_count_RNIQF5F5_4_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5831),
            .in3(N__10285),
            .lcout(\uu2.vbuf_tx_data_rdy ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI2U5E_10_LC_4_12_4 .C_ON=1'b0;
    defparam \uu2.l_count_RNI2U5E_10_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI2U5E_10_LC_4_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.l_count_RNI2U5E_10_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__5695),
            .in2(_gnd_net_),
            .in3(N__6064),
            .lcout(\uu2.un3_r_clk_en_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI89GK1_2_LC_4_12_5 .C_ON=1'b0;
    defparam \uu2.l_count_RNI89GK1_2_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI89GK1_2_LC_4_12_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uu2.l_count_RNI89GK1_2_LC_4_12_5  (
            .in0(N__6097),
            .in1(N__5768),
            .in2(N__6137),
            .in3(N__5742),
            .lcout(\uu2.un3_r_clk_en_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_7_LC_4_12_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_4_12_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_7_LC_4_12_6 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \buart.Z_tx.shifter_7_LC_4_12_6  (
            .in0(N__10287),
            .in1(N__5705),
            .in2(N__10508),
            .in3(N__7037),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13388),
            .ce(N__8588),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_8_LC_4_12_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_4_12_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_8_LC_4_12_7 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \buart.Z_tx.shifter_8_LC_4_12_7  (
            .in0(N__7262),
            .in1(N__10477),
            .in2(_gnd_net_),
            .in3(N__10288),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13388),
            .ce(N__8588),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_10__un372_ci_LC_4_13_0 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_10__un372_ci_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_10__un372_ci_LC_4_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_10__un372_ci_LC_4_13_0  (
            .in0(N__6036),
            .in1(N__6134),
            .in2(N__6151),
            .in3(N__6112),
            .lcout(),
            .ltout(\uu2.un372_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_10_LC_4_13_1 .C_ON=1'b0;
    defparam \uu2.l_count_10_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_10_LC_4_13_1 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \uu2.l_count_10_LC_4_13_1  (
            .in0(N__10469),
            .in1(_gnd_net_),
            .in2(N__5699),
            .in3(N__5696),
            .lcout(\uu2.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13384),
            .ce(),
            .sr(N__12301));
    defparam \uu2.l_count_8_LC_4_13_2 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_4_13_2 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_8_LC_4_13_2 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.l_count_8_LC_4_13_2  (
            .in0(N__6037),
            .in1(_gnd_net_),
            .in2(N__6152),
            .in3(N__6135),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13384),
            .ce(),
            .sr(N__12301));
    defparam \uu2.vbuf_count.counter_gen_label_10__un372_ci_8_1_LC_4_13_3 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_10__un372_ci_8_1_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_10__un372_ci_8_1_LC_4_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_10__un372_ci_8_1_LC_4_13_3  (
            .in0(N__6092),
            .in1(N__6173),
            .in2(N__6015),
            .in3(N__6065),
            .lcout(\uu2.vbuf_count.un372_ci_8_1 ),
            .ltout(\uu2.vbuf_count.un372_ci_8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_9_LC_4_13_4 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_4_13_4 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_9_LC_4_13_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.l_count_9_LC_4_13_4  (
            .in0(N__6039),
            .in1(N__6136),
            .in2(N__6116),
            .in3(N__6113),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13384),
            .ce(),
            .sr(N__12301));
    defparam \uu2.l_count_6_LC_4_13_5 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_4_13_5 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_6_LC_4_13_5 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.l_count_6_LC_4_13_5  (
            .in0(N__6093),
            .in1(N__6043),
            .in2(N__6017),
            .in3(N__6067),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13384),
            .ce(),
            .sr(N__12301));
    defparam \uu2.l_count_5_LC_4_13_6 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_4_13_6 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_5_LC_4_13_6 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu2.l_count_5_LC_4_13_6  (
            .in0(N__6066),
            .in1(N__6009),
            .in2(N__6044),
            .in3(N__10471),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13384),
            .ce(),
            .sr(N__12301));
    defparam \uu2.l_count_4_LC_4_13_7 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_4_13_7 .SEQ_MODE=4'b1000;
    defparam \uu2.l_count_4_LC_4_13_7 .LUT_INIT=16'b0001010000010100;
    LogicCell40 \uu2.l_count_4_LC_4_13_7  (
            .in0(N__10470),
            .in1(N__6038),
            .in2(N__6016),
            .in3(_gnd_net_),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13384),
            .ce(),
            .sr(N__12301));
    defparam \Lab_UT.secuu0.l_count_RNI24E71_11_LC_5_4_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNI24E71_11_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNI24E71_11_LC_5_4_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNI24E71_11_LC_5_4_0  (
            .in0(N__6254),
            .in1(N__6628),
            .in2(N__5978),
            .in3(N__6285),
            .lcout(\Lab_UT.secuu0.un4_l_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_RNI8TM21_5_LC_5_4_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNI8TM21_5_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNI8TM21_5_LC_5_4_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.secuu0.l_count_RNI8TM21_5_LC_5_4_4  (
            .in0(N__5953),
            .in1(N__5936),
            .in2(N__5912),
            .in3(N__6608),
            .lcout(),
            .ltout(\Lab_UT.secuu0.un4_l_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_RNI9GD02_18_LC_5_4_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNI9GD02_18_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNI9GD02_18_LC_5_4_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNI9GD02_18_LC_5_4_5  (
            .in0(N__6229),
            .in1(N__5892),
            .in2(N__5879),
            .in3(N__6517),
            .lcout(),
            .ltout(\Lab_UT.secuu0.un4_l_count_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_RNI82GM6_3_LC_5_4_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNI82GM6_3_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNI82GM6_3_LC_5_4_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNI82GM6_3_LC_5_4_6  (
            .in0(N__6353),
            .in1(N__6686),
            .in2(N__6347),
            .in3(N__6344),
            .lcout(\Lab_UT.secuu0.un4_l_count_0 ),
            .ltout(\Lab_UT.secuu0.un4_l_count_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.delay_line_RNILBAI7_1_LC_5_4_7 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.delay_line_RNILBAI7_1_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.delay_line_RNILBAI7_1_LC_5_4_7 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \Lab_UT.secuu0.delay_line_RNILBAI7_1_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(N__6335),
            .in2(N__6329),
            .in3(N__6325),
            .lcout(\Lab_UT.secuu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_0_LC_5_5_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_0_LC_5_5_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_0_LC_5_5_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.secuu0.l_count_0_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__6460),
            .in2(_gnd_net_),
            .in3(N__6634),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13423),
            .ce(N__6374),
            .sr(N__12312));
    defparam \Lab_UT.secuu0.l_count_11_LC_5_5_2 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_11_LC_5_5_2 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_11_LC_5_5_2 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Lab_UT.secuu0.l_count_11_LC_5_5_2  (
            .in0(N__6461),
            .in1(N__6577),
            .in2(N__6296),
            .in3(N__6287),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13423),
            .ce(N__6374),
            .sr(N__12312));
    defparam \Lab_UT.secuu0.l_count_16_LC_5_5_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_16_LC_5_5_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_16_LC_5_5_3 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \Lab_UT.secuu0.l_count_16_LC_5_5_3  (
            .in0(N__6267),
            .in1(N__6462),
            .in2(N__6584),
            .in3(N__6252),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13423),
            .ce(N__6374),
            .sr(N__12312));
    defparam \Lab_UT.secuu0.l_count_17_LC_5_5_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_17_LC_5_5_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_17_LC_5_5_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \Lab_UT.secuu0.l_count_17_LC_5_5_4  (
            .in0(N__6253),
            .in1(N__6268),
            .in2(N__6583),
            .in3(N__6187),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13423),
            .ce(N__6374),
            .sr(N__12312));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_18__un263_ci_LC_5_5_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_18__un263_ci_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_18__un263_ci_LC_5_5_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_18__un263_ci_LC_5_5_5  (
            .in0(N__6186),
            .in1(N__6568),
            .in2(N__6269),
            .in3(N__6251),
            .lcout(),
            .ltout(\Lab_UT.secuu0.un263_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_18_LC_5_5_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_18_LC_5_5_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_18_LC_5_5_6 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \Lab_UT.secuu0.l_count_18_LC_5_5_6  (
            .in0(N__6463),
            .in1(_gnd_net_),
            .in2(N__6233),
            .in3(N__6230),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13423),
            .ce(N__6374),
            .sr(N__12312));
    defparam \Lab_UT.secuu0.l_count_RNIRDS11_3_LC_5_5_7 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_RNIRDS11_3_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.l_count_RNIRDS11_3_LC_5_5_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.secuu0.l_count_RNIRDS11_3_LC_5_5_7  (
            .in0(N__6208),
            .in1(N__6666),
            .in2(N__6188),
            .in3(N__6390),
            .lcout(\Lab_UT.secuu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_3_LC_5_6_0 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_3_LC_5_6_0 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_3_LC_5_6_0 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \Lab_UT.secuu0.l_count_3_LC_5_6_0  (
            .in0(N__6668),
            .in1(N__6484),
            .in2(N__6680),
            .in3(N__6653),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13416),
            .ce(N__6373),
            .sr(N__12310));
    defparam \Lab_UT.secuu0.l_count_1_LC_5_6_1 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_1_LC_5_6_1 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_1_LC_5_6_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.secuu0.l_count_1_LC_5_6_1  (
            .in0(N__6607),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6633),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13416),
            .ce(N__6373),
            .sr(N__12310));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_1_LC_5_6_2 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_1_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_1_LC_5_6_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_1_LC_5_6_2  (
            .in0(N__6632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6606),
            .lcout(\Lab_UT.secuu0.un87_ci ),
            .ltout(\Lab_UT.secuu0.un87_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_2_LC_5_6_3 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_2_LC_5_6_3 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_2_LC_5_6_3 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \Lab_UT.secuu0.l_count_2_LC_5_6_3  (
            .in0(N__6652),
            .in1(_gnd_net_),
            .in2(N__6671),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13416),
            .ce(N__6373),
            .sr(N__12310));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_6_LC_5_6_4 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_6_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_6_LC_5_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_6_LC_5_6_4  (
            .in0(N__6667),
            .in1(N__6651),
            .in2(N__6635),
            .in3(N__6605),
            .lcout(\Lab_UT.secuu0.un109_ci ),
            .ltout(\Lab_UT.secuu0.un109_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_8_LC_5_6_5 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_8_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_8_LC_5_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.secuu0.vbuf_count_cntrl1.counter_gen_label_10__un175_ci_8_LC_5_6_5  (
            .in0(N__6529),
            .in1(N__6512),
            .in2(N__6587),
            .in3(N__6391),
            .lcout(\Lab_UT.secuu0.un153_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.l_count_6_LC_5_6_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_6_LC_5_6_6 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_6_LC_5_6_6 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \Lab_UT.secuu0.l_count_6_LC_5_6_6  (
            .in0(N__6513),
            .in1(N__6530),
            .in2(N__6421),
            .in3(N__6482),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13416),
            .ce(N__6373),
            .sr(N__12310));
    defparam \Lab_UT.secuu0.l_count_7_LC_5_6_7 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.l_count_7_LC_5_6_7 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.secuu0.l_count_7_LC_5_6_7 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \Lab_UT.secuu0.l_count_7_LC_5_6_7  (
            .in0(N__6483),
            .in1(N__6434),
            .in2(N__6395),
            .in3(N__6416),
            .lcout(\Lab_UT.secuu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13416),
            .ce(N__6373),
            .sr(N__12310));
    defparam \resetGen.reset_count_2_LC_5_7_0 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_5_7_0 .LUT_INIT=16'b0000000011100001;
    LogicCell40 \resetGen.reset_count_2_LC_5_7_0  (
            .in0(N__6809),
            .in1(N__6719),
            .in2(N__6776),
            .in3(N__6753),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13411),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_5_7_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_5_7_1 .LUT_INIT=16'b0100010001000001;
    LogicCell40 \resetGen.reset_count_3_LC_5_7_1  (
            .in0(N__6754),
            .in1(N__6739),
            .in2(N__6727),
            .in3(N__6761),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13411),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_5_7_2 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_5_7_2 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \resetGen.reset_count_0_LC_5_7_2  (
            .in0(N__6802),
            .in1(N__6717),
            .in2(_gnd_net_),
            .in3(N__6752),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13411),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.un3_reset_count_i_a3_LC_5_7_3 .C_ON=1'b0;
    defparam \resetGen.un3_reset_count_i_a3_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.un3_reset_count_i_a3_LC_5_7_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \resetGen.un3_reset_count_i_a3_LC_5_7_3  (
            .in0(N__13463),
            .in1(N__10724),
            .in2(N__12172),
            .in3(N__7565),
            .lcout(\resetGen.N_104 ),
            .ltout(\resetGen.N_104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_5_7_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_5_7_4 .LUT_INIT=16'b0000110100000010;
    LogicCell40 \resetGen.reset_count_1_LC_5_7_4  (
            .in0(N__6803),
            .in1(N__6718),
            .in2(N__6812),
            .in3(N__6788),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13411),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNO_0_2_LC_5_7_5 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_2_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_2_LC_5_7_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \resetGen.reset_count_RNO_0_2_LC_5_7_5  (
            .in0(N__6787),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6800),
            .lcout(\resetGen.N_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNITEEC1_2_LC_5_7_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNITEEC1_2_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNITEEC1_2_LC_5_7_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \resetGen.reset_count_RNITEEC1_2_LC_5_7_6  (
            .in0(N__6801),
            .in1(N__6786),
            .in2(_gnd_net_),
            .in3(N__6772),
            .lcout(\resetGen.N_86 ),
            .ltout(\resetGen.N_86_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_5_7_7 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_5_7_7 .LUT_INIT=16'b0101010100000100;
    LogicCell40 \resetGen.reset_count_4_LC_5_7_7  (
            .in0(N__6755),
            .in1(N__6740),
            .in2(N__6731),
            .in3(N__6723),
            .lcout(\resetGen.reset_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13411),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_5_8_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_5_8_0 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_44_LC_5_8_0  (
            .in0(N__11864),
            .in1(N__9704),
            .in2(N__9871),
            .in3(N__9965),
            .lcout(),
            .ltout(\uu2.mem0.g2_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_5_8_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_5_8_1 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_25_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__6845),
            .in2(N__6869),
            .in3(N__9440),
            .lcout(\uu2.mem0.g0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_5_8_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_5_8_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_40_LC_5_8_2  (
            .in0(N__9861),
            .in1(N__8473),
            .in2(_gnd_net_),
            .in3(N__8548),
            .lcout(),
            .ltout(\uu2.mem0.g0_i_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_5_8_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_5_8_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_24_LC_5_8_3  (
            .in0(N__7688),
            .in1(N__11865),
            .in2(N__6860),
            .in3(N__12682),
            .lcout(\uu2.mem0.w_data_displaying_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_5_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_5_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_52_LC_5_8_4  (
            .in0(N__9598),
            .in1(N__9540),
            .in2(N__9242),
            .in3(N__9162),
            .lcout(\uu2.mem0.g1_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_5_8_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_5_8_5 .LUT_INIT=16'b0010000000100101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_42_LC_5_8_5  (
            .in0(N__8547),
            .in1(N__12681),
            .in2(N__8477),
            .in3(N__12073),
            .lcout(\uu2.mem0.N_10_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_5_8_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_5_8_6 .LUT_INIT=16'b1100110011011110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_48_LC_5_8_6  (
            .in0(N__12072),
            .in1(N__9869),
            .in2(N__12698),
            .in3(N__8417),
            .lcout(\uu2.mem0.g1_1_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_5_8_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_5_8_7 .LUT_INIT=16'b1100001111100011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_32_LC_5_8_7  (
            .in0(N__10936),
            .in1(N__10697),
            .in2(N__10625),
            .in3(N__11416),
            .lcout(\uu2.mem0.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_5_9_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_5_9_0 .LUT_INIT=16'b0000001000000011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_27_LC_5_9_0  (
            .in0(N__8492),
            .in1(N__9705),
            .in2(N__6830),
            .in3(N__9964),
            .lcout(\uu2.mem0.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_5_9_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_5_9_1 .LUT_INIT=16'b0000000110101011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_60_LC_5_9_1  (
            .in0(N__12370),
            .in1(N__9074),
            .in2(N__9257),
            .in3(N__9235),
            .lcout(\uu2.mem0.g0_i_6_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_5_9_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_5_9_2 .LUT_INIT=16'b0111001001111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_38_LC_5_9_2  (
            .in0(N__9236),
            .in1(N__9062),
            .in2(N__7766),
            .in3(N__9164),
            .lcout(\uu2.mem0.g0_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_5_9_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_5_9_3 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_59_LC_5_9_3  (
            .in0(N__9800),
            .in1(N__9605),
            .in2(N__12371),
            .in3(N__9545),
            .lcout(),
            .ltout(\uu2.mem0.N_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_5_9_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_5_9_4 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_39_LC_5_9_4  (
            .in0(N__6899),
            .in1(N__8328),
            .in2(N__6893),
            .in3(N__9163),
            .lcout(\uu2.mem0.g0_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_5_9_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_5_9_5 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_53_LC_5_9_5  (
            .in0(N__11683),
            .in1(N__9422),
            .in2(N__9968),
            .in3(N__8546),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dicfsm.cState_LC_5_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrluu0.dicfsm.cState_LC_5_9_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \Lab_UT.dictrluu0.dicfsm.cState_LC_5_9_7  (
            .in0(N__10059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(Lab_UT_dicRun),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13399),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_5_10_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_5_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__6944),
            .in2(N__6926),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_5_10_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_5_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7160),
            .in3(N__6878),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_5_10_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_5_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_5_10_2  (
            .in0(N__7443),
            .in1(N__6992),
            .in2(_gnd_net_),
            .in3(N__6875),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__13394),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_5_10_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_5_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__6976),
            .in2(_gnd_net_),
            .in3(N__6872),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_5_10_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_5_10_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_5_10_4  (
            .in0(N__7445),
            .in1(N__7295),
            .in2(N__6962),
            .in3(N__7031),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13394),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNII0231_0_LC_5_10_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNII0231_0_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNII0231_0_LC_5_10_5 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNII0231_0_LC_5_10_5  (
            .in0(N__11794),
            .in1(N__7442),
            .in2(N__7300),
            .in3(N__7537),
            .lcout(\buart.Z_rx.bitcounte_0_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_10_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_10_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_5_10_6  (
            .in0(N__7444),
            .in1(N__7028),
            .in2(N__6980),
            .in3(N__7296),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13394),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_5_10_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_5_10_7 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_37_LC_5_10_7  (
            .in0(N__12694),
            .in1(N__8407),
            .in2(N__11244),
            .in3(N__8324),
            .lcout(\uu2.mem0.g0_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_5_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_5_11_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_5_11_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_5_11_0  (
            .in0(N__7454),
            .in1(N__6924),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13389),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_RNIVHME_0_LC_5_11_1 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNIVHME_0_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNIVHME_0_LC_5_11_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \buart.Z_rx.hh_RNIVHME_0_LC_5_11_1  (
            .in0(N__7858),
            .in1(N__7003),
            .in2(_gnd_net_),
            .in3(N__7538),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(\buart.Z_rx.startbit_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_5_11_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_5_11_2 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_5_11_2  (
            .in0(N__6943),
            .in1(_gnd_net_),
            .in2(N__7007),
            .in3(N__6925),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13389),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_1_LC_5_11_3 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.hh_1_LC_5_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7004),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13389),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_5_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_5_11_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_5_11_5  (
            .in0(N__6991),
            .in1(N__6975),
            .in2(N__6961),
            .in3(N__6942),
            .lcout(),
            .ltout(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_5_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_5_11_6 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__7155),
            .in2(N__6929),
            .in3(N__6923),
            .lcout(\buart.Z_rx.ser_clk ),
            .ltout(\buart.Z_rx.ser_clk_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_5_11_7 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_5_11_7 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_5_11_7  (
            .in0(N__7156),
            .in1(N__7453),
            .in2(N__7169),
            .in3(N__7166),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13389),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_esr_0_LC_5_12_0 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_0_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_0_LC_5_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_0_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7142),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13385),
            .ce(N__7253),
            .sr(N__12302));
    defparam \uu2.r_data_reg_esr_1_LC_5_12_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_1_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_1_LC_5_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_1_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7127),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13385),
            .ce(N__7253),
            .sr(N__12302));
    defparam \uu2.r_data_reg_esr_2_LC_5_12_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_2_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_2_LC_5_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_2_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7112),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13385),
            .ce(N__7253),
            .sr(N__12302));
    defparam \uu2.r_data_reg_esr_3_LC_5_12_3 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_3_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_3_LC_5_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_3_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7097),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13385),
            .ce(N__7253),
            .sr(N__12302));
    defparam \uu2.r_data_reg_esr_4_LC_5_12_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_4_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_4_LC_5_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_4_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7085),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13385),
            .ce(N__7253),
            .sr(N__12302));
    defparam \uu2.r_data_reg_esr_5_LC_5_12_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_5_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_5_LC_5_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_5_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7073),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13385),
            .ce(N__7253),
            .sr(N__12302));
    defparam \uu2.r_data_reg_esr_6_LC_5_12_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_6_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_6_LC_5_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_6_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7049),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13385),
            .ce(N__7253),
            .sr(N__12302));
    defparam \uu2.r_data_reg_esr_7_LC_5_12_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_esr_7_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_esr_7_LC_5_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_esr_7_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7274),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13385),
            .ce(N__7253),
            .sr(N__12302));
    defparam \buart.Z_tx.shifter_4_LC_5_13_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_4_LC_5_13_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \buart.Z_tx.shifter_4_LC_5_13_0  (
            .in0(N__10277),
            .in1(N__7235),
            .in2(N__7217),
            .in3(N__10488),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13381),
            .ce(N__8584),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_5_LC_5_13_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_5_LC_5_13_1 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \buart.Z_tx.shifter_5_LC_5_13_1  (
            .in0(N__7229),
            .in1(N__10485),
            .in2(N__10289),
            .in3(N__7223),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13381),
            .ce(N__8584),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_3_LC_5_13_2 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_3_LC_5_13_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \buart.Z_tx.shifter_3_LC_5_13_2  (
            .in0(N__10276),
            .in1(N__7208),
            .in2(N__7202),
            .in3(N__10487),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13381),
            .ce(N__8584),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_0_LC_5_13_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_0_LC_5_13_5 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \buart.Z_tx.shifter_0_LC_5_13_5  (
            .in0(N__7841),
            .in1(N__10484),
            .in2(_gnd_net_),
            .in3(N__10278),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13381),
            .ce(N__8584),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.uart_tx_LC_5_13_6 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.uart_tx_LC_5_13_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \buart.Z_tx.uart_tx_LC_5_13_6  (
            .in0(N__10275),
            .in1(N__7193),
            .in2(_gnd_net_),
            .in3(N__10486),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13381),
            .ce(N__8584),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_6_3_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_6_3_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_6_3_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_6_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_5_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__10754),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_5_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__7417),
            .in2(_gnd_net_),
            .in3(N__7172),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_5_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(N__10821),
            .in2(_gnd_net_),
            .in3(N__7346),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_5_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(N__10867),
            .in2(_gnd_net_),
            .in3(N__7343),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_4_LC_6_5_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_4_LC_6_5_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_e_0_4_LC_6_5_4 .LUT_INIT=16'b0001101101001110;
    LogicCell40 \buart.Z_rx.bitcount_e_0_4_LC_6_5_4  (
            .in0(N__7517),
            .in1(N__7557),
            .in2(N__7478),
            .in3(N__7340),
            .lcout(\buart.Z_rx.bitcountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13414),
            .ce(N__7391),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_0_LC_6_6_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_0_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_e_0_0_LC_6_6_1 .LUT_INIT=16'b0001001011011110;
    LogicCell40 \buart.Z_rx.bitcount_e_0_0_LC_6_6_1  (
            .in0(N__10761),
            .in1(N__7511),
            .in2(N__8892),
            .in3(N__7469),
            .lcout(buart__rx_bitcount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13409),
            .ce(N__7390),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_3_LC_6_6_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_3_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_e_0_3_LC_6_6_2 .LUT_INIT=16'b0101010100111100;
    LogicCell40 \buart.Z_rx.bitcount_e_0_3_LC_6_6_2  (
            .in0(N__7468),
            .in1(N__10868),
            .in2(N__7337),
            .in3(N__7513),
            .lcout(buart__rx_bitcount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13409),
            .ce(N__7390),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_2_LC_6_6_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_2_LC_6_6_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_e_0_2_LC_6_6_3 .LUT_INIT=16'b0001001011011110;
    LogicCell40 \buart.Z_rx.bitcount_e_0_2_LC_6_6_3  (
            .in0(N__10825),
            .in1(N__7512),
            .in2(N__7325),
            .in3(N__7470),
            .lcout(buart__rx_bitcount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13409),
            .ce(N__7390),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_6_6_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_6_6_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_15_LC_6_6_5  (
            .in0(N__9035),
            .in1(N__11242),
            .in2(_gnd_net_),
            .in3(N__11984),
            .lcout(\uu2.mem0.w_data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNI2B26_4_LC_6_7_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNI2B26_4_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNI2B26_4_LC_6_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNI2B26_4_LC_6_7_0  (
            .in0(N__10863),
            .in1(N__7559),
            .in2(N__7418),
            .in3(N__10819),
            .lcout(),
            .ltout(\buart.Z_rx.N_103_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNIBJOC_0_LC_6_7_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNIBJOC_0_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNIBJOC_0_LC_6_7_1 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNIBJOC_0_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(N__7304),
            .in2(N__7277),
            .in3(N__10753),
            .lcout(\buart.Z_rx.N_57_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_0_LC_6_7_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_0_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_0_LC_6_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNI8RI7_0_0_LC_6_7_2  (
            .in0(N__10783),
            .in1(N__10760),
            .in2(N__10872),
            .in3(N__10818),
            .lcout(bu_rx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.un3_reset_count_i_a3_7_LC_6_7_3 .C_ON=1'b0;
    defparam \resetGen.un3_reset_count_i_a3_7_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.un3_reset_count_i_a3_7_LC_6_7_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \resetGen.un3_reset_count_i_a3_7_LC_6_7_3  (
            .in0(N__10820),
            .in1(N__12218),
            .in2(N__10873),
            .in3(N__10782),
            .lcout(\resetGen.un3_reset_count_i_a3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNIH513_4_LC_6_7_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNIH513_4_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNIH513_4_LC_6_7_4 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNIH513_4_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(N__7558),
            .in2(_gnd_net_),
            .in3(N__7409),
            .lcout(N_87),
            .ltout(N_87_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_LC_6_7_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNI8RI7_0_LC_6_7_5 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNI8RI7_0_LC_6_7_5  (
            .in0(N__10817),
            .in1(N__10859),
            .in2(N__7541),
            .in3(N__10752),
            .lcout(\buart.Z_rx.N_91 ),
            .ltout(\buart.Z_rx.N_91_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_RNIGM5F_0_LC_6_7_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_RNIGM5F_0_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_e_0_RNIGM5F_0_LC_6_7_6 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \buart.Z_rx.bitcount_e_0_RNIGM5F_0_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7520),
            .in3(N__11781),
            .lcout(\buart.Z_rx.N_29_0_i_2 ),
            .ltout(\buart.Z_rx.N_29_0_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_e_0_1_LC_6_7_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_e_0_1_LC_6_7_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.bitcount_e_0_1_LC_6_7_7 .LUT_INIT=16'b0000011011110110;
    LogicCell40 \buart.Z_rx.bitcount_e_0_1_LC_6_7_7  (
            .in0(N__7410),
            .in1(N__7493),
            .in2(N__7481),
            .in3(N__7474),
            .lcout(\buart.Z_rx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13403),
            .ce(N__7383),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIAPHB1_5_LC_6_8_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIAPHB1_5_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIAPHB1_5_LC_6_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIAPHB1_5_LC_6_8_0  (
            .in0(N__11848),
            .in1(N__12683),
            .in2(N__9872),
            .in3(N__12059),
            .lcout(\uu2.Z_decfrac105_7_3 ),
            .ltout(\uu2.Z_decfrac105_7_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_8_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_8_1 .LUT_INIT=16'b0010000011101100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_6_8_1  (
            .in0(N__9371),
            .in1(N__11220),
            .in2(N__7358),
            .in3(N__10712),
            .lcout(\uu2.mem0.w_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_6_8_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_6_8_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_17_LC_6_8_2  (
            .in0(_gnd_net_),
            .in1(N__7657),
            .in2(_gnd_net_),
            .in3(N__9369),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_6_8_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_6_8_3 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_6_8_3  (
            .in0(N__11219),
            .in1(N__7706),
            .in2(N__7670),
            .in3(N__8230),
            .lcout(\uu2.mem0.w_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_6_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_6_8_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_18_LC_6_8_4  (
            .in0(N__12586),
            .in1(N__7658),
            .in2(_gnd_net_),
            .in3(N__9370),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_6_8_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_6_8_5 .LUT_INIT=16'b1101110111011000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_6_8_5  (
            .in0(N__11218),
            .in1(N__7697),
            .in2(N__7649),
            .in3(N__8231),
            .lcout(\uu2.mem0.w_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_5_LC_6_8_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_LC_6_8_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_LC_6_8_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_5_LC_6_8_6  (
            .in0(N__12497),
            .in1(N__12792),
            .in2(N__11863),
            .in3(N__12685),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_5C_net ),
            .ce(),
            .sr(N__12281));
    defparam \uu2.w_addr_displaying_4_LC_6_8_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_LC_6_8_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.w_addr_displaying_4_LC_6_8_7  (
            .in0(N__12684),
            .in1(N__12791),
            .in2(_gnd_net_),
            .in3(N__12498),
            .lcout(\uu2.w_addr_displayingZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_5C_net ),
            .ce(),
            .sr(N__12281));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_6_9_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_6_9_0 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_6_9_0  (
            .in0(N__9280),
            .in1(N__11102),
            .in2(N__7622),
            .in3(N__11030),
            .lcout(\uu2.mem0.w_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_0_LC_6_9_1 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_0_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_0_LC_6_9_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.un1_w_user_cr_0_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__8963),
            .in2(_gnd_net_),
            .in3(N__9320),
            .lcout(\uu2.un1_w_user_cr_0_0 ),
            .ltout(\uu2.un1_w_user_cr_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_wr_en_0_i_LC_6_9_2 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_6_9_2 .LUT_INIT=16'b0101110111011101;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_6_9_2  (
            .in0(N__7609),
            .in1(N__9279),
            .in2(N__7595),
            .in3(N__11101),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.rdy_LC_6_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.rdy_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.rdy_LC_6_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dspStr.rdy_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10154),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13392),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_6_9_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_6_9_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_34_LC_6_9_4  (
            .in0(N__8180),
            .in1(N__8207),
            .in2(N__7745),
            .in3(N__7772),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_6_9_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_6_9_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_20_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__9083),
            .in2(N__7730),
            .in3(N__7712),
            .lcout(),
            .ltout(\uu2.mem0.un1_segment3_m6_0_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_6_9_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_6_9_6 .LUT_INIT=16'b0111011001100110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_6_9_6  (
            .in0(N__11243),
            .in1(N__8216),
            .in2(N__7727),
            .in3(N__7676),
            .lcout(\uu2.mem0.w_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_6_9_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_6_9_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_35_LC_6_9_7  (
            .in0(N__8206),
            .in1(N__8179),
            .in2(_gnd_net_),
            .in3(N__7741),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_6_10_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_6_10_0 .LUT_INIT=16'b0110001001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_21_LC_6_10_0  (
            .in0(N__10695),
            .in1(N__10617),
            .in2(N__11945),
            .in3(N__10943),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_6_10_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_6_10_1 .LUT_INIT=16'b1110101011001010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_22_LC_6_10_1  (
            .in0(N__10942),
            .in1(N__10696),
            .in2(N__10624),
            .in3(N__11462),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_rep1_RNI56RN_LC_6_10_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_RNI56RN_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_0_rep1_RNI56RN_LC_6_10_2 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_RNI56RN_LC_6_10_2  (
            .in0(N__9410),
            .in1(N__8311),
            .in2(_gnd_net_),
            .in3(N__8520),
            .lcout(\uu2.g0_1_a5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_6_10_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_6_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_41_LC_6_10_3  (
            .in0(N__8312),
            .in1(N__11564),
            .in2(N__12078),
            .in3(N__8406),
            .lcout(\uu2.mem0.g0_i_a2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_6_10_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_6_10_4 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_16_LC_6_10_4  (
            .in0(N__7757),
            .in1(N__9467),
            .in2(N__8264),
            .in3(N__8339),
            .lcout(\uu2.mem0.N_8_tz_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.g0_LC_6_10_5 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.g0_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.g0_LC_6_10_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didpuu0.g0_LC_6_10_5  (
            .in0(N__13140),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13160),
            .lcout(),
            .ltout(led_c_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_6_10_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_6_10_6 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_56_LC_6_10_6  (
            .in0(N__9980),
            .in1(N__9699),
            .in2(N__7775),
            .in3(N__8429),
            .lcout(\uu2.mem0.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_6_10_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_6_10_7 .LUT_INIT=16'b0111111101000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_58_LC_6_10_7  (
            .in0(N__9419),
            .in1(N__13161),
            .in2(N__13145),
            .in3(N__9148),
            .lcout(\uu2.mem0.g0_i_5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_6_11_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_6_11_0 .LUT_INIT=16'b0100100000010010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_30_LC_6_11_0  (
            .in0(N__8397),
            .in1(N__12693),
            .in2(N__9703),
            .in3(N__12065),
            .lcout(\uu2.mem0.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_rep1_8_LC_6_11_1 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_rep1_8_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_rep1_8_LC_6_11_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_rep1_8_LC_6_11_1  (
            .in0(N__12798),
            .in1(N__9688),
            .in2(N__9763),
            .in3(N__8398),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_4_rep1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_8_rep1_LC_6_11_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_rep1_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_rep1_LC_6_11_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \uu2.w_addr_displaying_8_rep1_LC_6_11_2  (
            .in0(N__12500),
            .in1(_gnd_net_),
            .in2(N__7751),
            .in3(N__8408),
            .lcout(\uu2.w_addr_displaying_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8_rep1C_net ),
            .ce(),
            .sr(N__12285));
    defparam \uu2.w_addr_displaying_8_rep1_RNIN6OC_LC_6_11_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_rep1_RNIN6OC_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_8_rep1_RNIN6OC_LC_6_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_displaying_8_rep1_RNIN6OC_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(N__8309),
            .in2(_gnd_net_),
            .in3(N__8396),
            .lcout(),
            .ltout(\uu2.N_42_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI8V6F2_3_LC_6_11_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8V6F2_3_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8V6F2_3_LC_6_11_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI8V6F2_3_LC_6_11_4  (
            .in0(N__8594),
            .in1(N__12692),
            .in2(N__7748),
            .in3(N__12064),
            .lcout(\uu2.N_1482_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_7_rep1_LC_6_11_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_rep1_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_rep1_LC_6_11_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_7_rep1_LC_6_11_5  (
            .in0(N__12802),
            .in1(N__12499),
            .in2(N__9764),
            .in3(N__8310),
            .lcout(\uu2.w_addr_displaying_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8_rep1C_net ),
            .ce(),
            .sr(N__12285));
    defparam \uu2.w_addr_displaying_4_rep1_RNI65VM_LC_6_11_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep1_RNI65VM_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_4_rep1_RNI65VM_LC_6_11_6 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \uu2.w_addr_displaying_4_rep1_RNI65VM_LC_6_11_6  (
            .in0(N__8308),
            .in1(N__9132),
            .in2(N__8409),
            .in3(N__9204),
            .lcout(\uu2.g0_1_a5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_rep1_LC_6_11_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_rep1_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_rep1_LC_6_11_7 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \uu2.w_addr_displaying_4_rep1_LC_6_11_7  (
            .in0(N__9205),
            .in1(_gnd_net_),
            .in2(N__12808),
            .in3(N__12501),
            .lcout(\uu2.w_addr_displaying_4_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8_rep1C_net ),
            .ce(),
            .sr(N__12285));
    defparam \buart.Z_rx.shifter_7_LC_6_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_6_12_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_7_LC_6_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_LC_6_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7859),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13380),
            .ce(N__13255),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_6_13_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_6_13_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_1_LC_6_13_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \buart.Z_tx.shifter_1_LC_6_13_0  (
            .in0(N__7847),
            .in1(N__10517),
            .in2(N__7820),
            .in3(N__10279),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13378),
            .ce(N__8583),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_2_LC_6_13_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.shifter_2_LC_6_13_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \buart.Z_tx.shifter_2_LC_6_13_4  (
            .in0(N__7835),
            .in1(N__10518),
            .in2(N__7829),
            .in3(N__10280),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13378),
            .ce(N__8583),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un415_ci_LC_7_5_0 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un415_ci_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un415_ci_LC_7_5_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_4__un415_ci_LC_7_5_0  (
            .in0(N__7927),
            .in1(N__8110),
            .in2(N__7803),
            .in3(N__11277),
            .lcout(\uu2.un415_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_2_LC_7_5_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_2_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_2_LC_7_5_1 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_user_2_LC_7_5_1  (
            .in0(N__11280),
            .in1(N__7930),
            .in2(N__8119),
            .in3(N__8847),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__8777));
    defparam \uu2.vbuf_w_addr_user.result_1_3_LC_7_5_2 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.result_1_3_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.result_1_3_LC_7_5_2 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.vbuf_w_addr_user.result_1_3_LC_7_5_2  (
            .in0(N__7928),
            .in1(N__8111),
            .in2(N__7804),
            .in3(N__11278),
            .lcout(),
            .ltout(\uu2.o_adder_vbuf_w_addr_user_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_3_LC_7_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_3_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_3_LC_7_5_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \uu2.w_addr_user_3_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(N__7799),
            .in2(N__7811),
            .in3(N__8846),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__8777));
    defparam \uu2.w_addr_user_RNIDD1A_5_LC_7_5_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIDD1A_5_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIDD1A_5_LC_7_5_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_RNIDD1A_5_LC_7_5_6  (
            .in0(N__7792),
            .in1(N__7923),
            .in2(N__8032),
            .in3(N__11276),
            .lcout(\uu2.un2_w_addr_user_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_userZ0Z_1_LC_7_5_7 .C_ON=1'b0;
    defparam \uu2.w_addr_userZ0Z_1_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_userZ0Z_1_LC_7_5_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.w_addr_userZ0Z_1_LC_7_5_7  (
            .in0(N__11279),
            .in1(N__7929),
            .in2(_gnd_net_),
            .in3(N__8845),
            .lcout(\uu2.w_addr_userZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__8777));
    defparam \uu2.vbuf_w_addr_user.result_1_7_LC_7_6_0 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.result_1_7_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.result_1_7_LC_7_6_0 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.vbuf_w_addr_user.result_1_7_LC_7_6_0  (
            .in0(N__8140),
            .in1(N__7876),
            .in2(N__8085),
            .in3(N__7985),
            .lcout(),
            .ltout(\uu2.o_adder_vbuf_w_addr_user_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_7_LC_7_6_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_7_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_7_LC_7_6_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \uu2.w_addr_user_7_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__8141),
            .in2(N__7901),
            .in3(N__8842),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_7C_net ),
            .ce(),
            .sr(N__8786));
    defparam \uu2.w_addr_user_6_LC_7_6_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_6_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_6_LC_7_6_2 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_user_6_LC_7_6_2  (
            .in0(N__8844),
            .in1(N__7877),
            .in2(N__8086),
            .in3(N__7987),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_7C_net ),
            .ce(),
            .sr(N__8786));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_6_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_6_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_7_6_4  (
            .in0(N__8138),
            .in1(N__11217),
            .in2(_gnd_net_),
            .in3(N__9706),
            .lcout(\uu2.mem0.w_addr_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un459_ci_0_LC_7_6_5 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un459_ci_0_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un459_ci_0_LC_7_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_8__un459_ci_0_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(N__8074),
            .in2(_gnd_net_),
            .in3(N__8139),
            .lcout(),
            .ltout(\uu2.vbuf_w_addr_user.un459_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.result_1_8_LC_7_6_6 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.result_1_8_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.result_1_8_LC_7_6_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.vbuf_w_addr_user.result_1_8_LC_7_6_6  (
            .in0(N__7875),
            .in1(N__7986),
            .in2(N__7883),
            .in3(N__8165),
            .lcout(),
            .ltout(\uu2.o_adder_vbuf_w_addr_user_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_8_LC_7_6_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_8_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_8_LC_7_6_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uu2.w_addr_user_8_LC_7_6_7  (
            .in0(N__8166),
            .in1(_gnd_net_),
            .in2(N__7880),
            .in3(N__8843),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_7C_net ),
            .ce(),
            .sr(N__8786));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un437_ci_3_LC_7_7_0 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un437_ci_3_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un437_ci_3_LC_7_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_6__un437_ci_3_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__7968),
            .in2(_gnd_net_),
            .in3(N__8021),
            .lcout(\uu2.un437_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIKCH7_8_LC_7_7_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIKCH7_8_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIKCH7_8_LC_7_7_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uu2.w_addr_user_RNIKCH7_8_LC_7_7_1  (
            .in0(N__8167),
            .in1(N__8137),
            .in2(_gnd_net_),
            .in3(N__8115),
            .lcout(),
            .ltout(\uu2.un2_w_addr_user_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIDMJM_4_LC_7_7_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIDMJM_4_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIDMJM_4_LC_7_7_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu2.w_addr_user_RNIDMJM_4_LC_7_7_2  (
            .in0(N__8081),
            .in1(N__7966),
            .in2(N__8048),
            .in3(N__8045),
            .lcout(\uu2.un2_w_addr_user ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_7__un448_ci_5_LC_7_7_3 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_7__un448_ci_5_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_7__un448_ci_5_LC_7_7_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.vbuf_w_addr_displaying.counter_gen_label_7__un448_ci_5_LC_7_7_3  (
            .in0(N__9237),
            .in1(N__9582),
            .in2(_gnd_net_),
            .in3(N__9527),
            .lcout(\uu2.un448_ci_5 ),
            .ltout(\uu2.un448_ci_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_8_rep1_RNI5LHP1_LC_7_7_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_rep1_RNI5LHP1_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_8_rep1_RNI5LHP1_LC_7_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_8_rep1_RNI5LHP1_LC_7_7_4  (
            .in0(N__9463),
            .in1(N__8416),
            .in2(N__8036),
            .in3(N__8332),
            .lcout(\uu2.Z_decfrac106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_5_LC_7_7_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_5_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_5_LC_7_7_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_user_5_LC_7_7_5  (
            .in0(N__8855),
            .in1(N__7997),
            .in2(N__8031),
            .in3(N__7970),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__8781));
    defparam \uu2.w_addr_user_4_LC_7_7_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_4_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_4_LC_7_7_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.w_addr_user_4_LC_7_7_6  (
            .in0(N__7996),
            .in1(N__7969),
            .in2(_gnd_net_),
            .in3(N__8854),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__8781));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_7_7_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_7_7_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_7_7_7  (
            .in0(N__7967),
            .in1(N__11201),
            .in2(_gnd_net_),
            .in3(N__12686),
            .lcout(\uu2.mem0.w_addr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_64_LC_7_8_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_64_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_64_LC_7_8_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_64_LC_7_8_0  (
            .in0(_gnd_net_),
            .in1(N__9523),
            .in2(_gnd_net_),
            .in3(N__9155),
            .lcout(),
            .ltout(\uu2.mem0.g0_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_7_8_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_7_8_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_46_LC_7_8_1  (
            .in0(N__12676),
            .in1(N__9870),
            .in2(N__7937),
            .in3(N__9361),
            .lcout(),
            .ltout(\uu2.mem0.w_data_ns_1_1_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_7_8_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_7_8_2 .LUT_INIT=16'b0111011101000111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_26_LC_7_8_2  (
            .in0(N__8741),
            .in1(N__11183),
            .in2(N__8234),
            .in3(N__8229),
            .lcout(\uu2.mem0.w_data_ns_1_0_0_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_5_rep1_LC_7_8_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_rep1_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_rep1_LC_7_8_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_5_rep1_LC_7_8_3  (
            .in0(N__12677),
            .in1(N__12759),
            .in2(N__9539),
            .in3(N__12467),
            .lcout(\uu2.w_addr_displaying_5_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_5_rep1C_net ),
            .ce(),
            .sr(N__12282));
    defparam \uu2.w_addr_displaying_6_rep1_RNI6D891_LC_7_8_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_rep1_RNI6D891_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_6_rep1_RNI6D891_LC_7_8_4 .LUT_INIT=16'b0000011111111111;
    LogicCell40 \uu2.w_addr_displaying_6_rep1_RNI6D891_LC_7_8_4  (
            .in0(N__9581),
            .in1(N__9522),
            .in2(N__12705),
            .in3(N__12049),
            .lcout(),
            .ltout(\uu2.g0_1_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIRTT92_8_LC_7_8_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIRTT92_8_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIRTT92_8_LC_7_8_5 .LUT_INIT=16'b0000010100010111;
    LogicCell40 \uu2.w_addr_displaying_RNIRTT92_8_LC_7_8_5  (
            .in0(N__12675),
            .in1(N__9695),
            .in2(N__8210),
            .in3(N__9957),
            .lcout(\uu2.g0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_LC_7_8_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_LC_7_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.w_addr_displaying_3_LC_7_8_6  (
            .in0(N__11999),
            .in1(N__12465),
            .in2(_gnd_net_),
            .in3(N__12050),
            .lcout(\uu2.w_addr_displayingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_5_rep1C_net ),
            .ce(),
            .sr(N__12282));
    defparam \uu2.w_addr_displaying_6_rep1_LC_7_8_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_rep1_LC_7_8_7 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_6_rep1_LC_7_8_7 .LUT_INIT=16'b1101111010101010;
    LogicCell40 \uu2.w_addr_displaying_6_rep1_LC_7_8_7  (
            .in0(N__9589),
            .in1(N__9901),
            .in2(N__11825),
            .in3(N__12468),
            .lcout(\uu2.w_addr_displaying_6_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_5_rep1C_net ),
            .ce(),
            .sr(N__12282));
    defparam \uu2.w_addr_displaying_RNI2AJ42_5_LC_7_9_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI2AJ42_5_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI2AJ42_5_LC_7_9_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \uu2.w_addr_displaying_RNI2AJ42_5_LC_7_9_2  (
            .in0(N__9843),
            .in1(N__11847),
            .in2(N__8198),
            .in3(N__8189),
            .lcout(\uu2.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_rep1_LC_7_9_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_rep1_LC_7_9_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_LC_7_9_4  (
            .in0(N__12462),
            .in1(N__11677),
            .in2(N__12601),
            .in3(N__9420),
            .lcout(\uu2.w_addr_displaying_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__12284));
    defparam \uu2.w_addr_displaying_2_LC_7_9_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_7_9_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_2_LC_7_9_5  (
            .in0(N__11676),
            .in1(N__12591),
            .in2(N__11592),
            .in3(N__12464),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__12284));
    defparam \uu2.w_addr_displaying_RNIUCHB1_2_LC_7_9_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIUCHB1_2_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIUCHB1_2_LC_7_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIUCHB1_2_LC_7_9_6  (
            .in0(N__11571),
            .in1(N__11674),
            .in2(N__12600),
            .in3(N__12063),
            .lcout(\uu2.un15_w_data_displaying_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_LC_7_9_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_LC_7_9_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.w_addr_displaying_1_LC_7_9_7  (
            .in0(N__11675),
            .in1(N__12590),
            .in2(_gnd_net_),
            .in3(N__12463),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__12284));
    defparam \uu2.w_addr_displaying_6_rep1_RNIAP701_LC_7_10_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_rep1_RNIAP701_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_6_rep1_RNIAP701_LC_7_10_0 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \uu2.w_addr_displaying_6_rep1_RNIAP701_LC_7_10_0  (
            .in0(N__8313),
            .in1(N__8399),
            .in2(N__9544),
            .in3(N__9603),
            .lcout(\uu2.g1_0_1 ),
            .ltout(\uu2.g1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_7_10_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_7_10_1 .LUT_INIT=16'b1111100110011001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_50_LC_7_10_1  (
            .in0(N__9210),
            .in1(N__9135),
            .in2(N__8351),
            .in3(N__8251),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_7_10_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_7_10_2 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_28_LC_7_10_2  (
            .in0(N__8252),
            .in1(N__8240),
            .in2(N__8348),
            .in3(N__8345),
            .lcout(\uu2.mem0.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_7_10_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_7_10_3 .LUT_INIT=16'b1111100100001001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_51_LC_7_10_3  (
            .in0(N__9209),
            .in1(N__9134),
            .in2(N__9966),
            .in3(N__8250),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_7_10_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_7_10_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_29_LC_7_10_4  (
            .in0(N__8314),
            .in1(_gnd_net_),
            .in2(N__8267),
            .in3(N__9604),
            .lcout(\uu2.mem0.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI7RCN_4_LC_7_10_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI7RCN_4_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI7RCN_4_LC_7_10_5 .LUT_INIT=16'b0000101000010001;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI7RCN_4_LC_7_10_5  (
            .in0(N__8521),
            .in1(N__9133),
            .in2(N__10019),
            .in3(N__8461),
            .lcout(\uu2.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_7_10_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_7_10_6 .LUT_INIT=16'b0100100000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_49_LC_7_10_6  (
            .in0(N__8462),
            .in1(N__9534),
            .in2(N__9421),
            .in3(N__9602),
            .lcout(\uu2.mem0.g1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_rep1_LC_7_10_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_rep1_LC_7_10_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_LC_7_10_7  (
            .in0(N__12493),
            .in1(_gnd_net_),
            .in2(N__8534),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displaying_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0_rep1C_net ),
            .ce(),
            .sr(N__12286));
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_7_11_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_7_11_0 .LUT_INIT=16'b0000110000010001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_47_LC_7_11_0  (
            .in0(N__9136),
            .in1(N__8466),
            .in2(N__9228),
            .in3(N__8525),
            .lcout(\uu2.mem0.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_rep1_3_LC_7_11_1 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_rep1_3_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_rep1_3_LC_7_11_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_rep1_3_LC_7_11_1  (
            .in0(N__11586),
            .in1(N__11692),
            .in2(N__12602),
            .in3(N__9137),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_4_rep1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_rep1_LC_7_11_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_rep1_LC_7_11_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_LC_7_11_2  (
            .in0(N__9138),
            .in1(_gnd_net_),
            .in2(N__8480),
            .in3(N__12502),
            .lcout(\uu2.w_addr_displaying_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__12288));
    defparam \uu2.w_addr_displaying_1_rep1_LC_7_11_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_rep1_LC_7_11_3 .LUT_INIT=16'b0110101001101010;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_LC_7_11_3  (
            .in0(N__8467),
            .in1(N__12599),
            .in2(N__12509),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displaying_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__12288));
    defparam \uu2.w_addr_displaying_fast_2_LC_7_11_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_2_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_2_LC_7_11_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_fast_2_LC_7_11_4  (
            .in0(N__11693),
            .in1(N__12504),
            .in2(N__8441),
            .in3(N__12598),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__12288));
    defparam \uu2.mem0.ram512X8_inst_RNO_66_LC_7_11_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_66_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_66_LC_7_11_5 .LUT_INIT=16'b1101010110101111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_66_LC_7_11_5  (
            .in0(N__11633),
            .in1(N__8423),
            .in2(N__10018),
            .in3(N__8437),
            .lcout(\uu2.mem0.un1_segment4_0_i_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_4_LC_7_11_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_4_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_4_LC_7_11_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.w_addr_displaying_fast_4_LC_7_11_6  (
            .in0(N__10014),
            .in1(N__12503),
            .in2(_gnd_net_),
            .in3(N__12803),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__12288));
    defparam \uu2.mem0.ram512X8_inst_RNO_71_LC_7_12_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_71_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_71_LC_7_12_0 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_71_LC_7_12_0  (
            .in0(N__13030),
            .in1(N__12860),
            .in2(N__12983),
            .in3(N__13209),
            .lcout(\uu2.mem0.un1_segment4_0_i_i_a5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_RNIUTLC1_2_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_RNIUTLC1_2_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpsones.q_RNIUTLC1_2_LC_7_12_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_RNIUTLC1_2_LC_7_12_1  (
            .in0(N__13210),
            .in1(N__13032),
            .in2(N__12876),
            .in3(N__12966),
            .lcout(\Lab_UT.didpuu0.didpsones.q13_0 ),
            .ltout(\Lab_UT.didpuu0.didpsones.q13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_2_LC_7_12_2 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_2_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpsones.q_2_LC_7_12_2 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_2_LC_7_12_2  (
            .in0(N__10124),
            .in1(N__11732),
            .in2(N__8597),
            .in3(N__10076),
            .lcout(Lab_UT_di_Sones_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13386),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.g0_3_0_LC_7_12_7 .C_ON=1'b0;
    defparam \uu2.g0_3_0_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \uu2.g0_3_0_LC_7_12_7 .LUT_INIT=16'b1111011001111101;
    LogicCell40 \uu2.g0_3_0_LC_7_12_7  (
            .in0(N__13208),
            .in1(N__12962),
            .in2(N__12875),
            .in3(N__13031),
            .lcout(\uu2.g0_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_7_13_0 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_7_13_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_7_13_0  (
            .in0(N__8639),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8659),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13382),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_7_13_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_7_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8638),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13382),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_RNO_LC_7_13_3 .C_ON=1'b0;
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_RNO_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_RNO_LC_7_13_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \buart.Z_tx.un1_bitcount_cry_0_c_RNO_LC_7_13_3  (
            .in0(N__10236),
            .in1(N__10372),
            .in2(_gnd_net_),
            .in3(N__10317),
            .lcout(\buart.Z_tx.un1_bitcount_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIV5CT5_1_LC_7_13_4 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIV5CT5_1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIV5CT5_1_LC_7_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIV5CT5_1_LC_7_13_4  (
            .in0(N__10318),
            .in1(N__10509),
            .in2(_gnd_net_),
            .in3(N__10237),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_1_LC_7_13_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_1_LC_7_13_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_7_13_6  (
            .in0(N__10516),
            .in1(N__10239),
            .in2(_gnd_net_),
            .in3(N__10028),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13382),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_0_LC_7_13_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_0_LC_7_13_7 .LUT_INIT=16'b0001100101001100;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_7_13_7  (
            .in0(N__10238),
            .in1(N__10371),
            .in2(N__10519),
            .in3(N__10319),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13382),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_7_14_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_7_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__8637),
            .in2(N__8660),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_7_14_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_7_14_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8618),
            .in3(N__8723),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__13379),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_7_14_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_7_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_7_14_2  (
            .in0(N__10324),
            .in1(N__8669),
            .in2(_gnd_net_),
            .in3(N__8720),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__13379),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_7_14_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_7_14_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8696),
            .in3(N__8717),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__13379),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_7_14_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_7_14_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_7_14_4  (
            .in0(N__10325),
            .in1(_gnd_net_),
            .in2(N__8708),
            .in3(N__8714),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__13379),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_7_14_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_7_14_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_7_14_5  (
            .in0(N__8683),
            .in1(N__10323),
            .in2(_gnd_net_),
            .in3(N__8711),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13379),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_7_14_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_7_14_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_7_14_6  (
            .in0(N__8704),
            .in1(N__8692),
            .in2(N__8684),
            .in3(N__8668),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_7_14_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_7_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_7_14_7  (
            .in0(N__8655),
            .in1(N__8636),
            .in2(N__8617),
            .in3(N__8603),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_0_LC_8_4_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_0_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_0_LC_8_4_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_user_0_LC_8_4_0  (
            .in0(_gnd_net_),
            .in1(N__11284),
            .in2(_gnd_net_),
            .in3(N__8853),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_0C_net ),
            .ce(),
            .sr(N__8785));
    defparam \uu2.w_addr_user_2_1_LC_8_5_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_2_1_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_2_1_LC_8_5_0 .LUT_INIT=16'b0000111100001011;
    LogicCell40 \uu2.w_addr_user_2_1_LC_8_5_0  (
            .in0(N__11905),
            .in1(N__8942),
            .in2(N__10691),
            .in3(N__11982),
            .lcout(),
            .ltout(\uu2.w_addr_user_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNILAII7_4_LC_8_5_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNILAII7_4_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNILAII7_4_LC_8_5_1 .LUT_INIT=16'b1110111111101110;
    LogicCell40 \uu2.w_addr_user_RNILAII7_4_LC_8_5_1  (
            .in0(N__8921),
            .in1(N__10065),
            .in2(N__8792),
            .in3(N__11095),
            .lcout(),
            .ltout(\uu2.w_addr_userZ2Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIT1MGD_4_LC_8_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIT1MGD_4_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIT1MGD_4_LC_8_5_2 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \uu2.w_addr_user_RNIT1MGD_4_LC_8_5_2  (
            .in0(N__8750),
            .in1(N__8927),
            .in2(N__8789),
            .in3(N__8807),
            .lcout(\uu2.w_addr_user_RNIT1MGDZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_1_LC_8_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_1_LC_8_5_3 .LUT_INIT=16'b0001111100001010;
    LogicCell40 \uu2.w_addr_user_1_LC_8_5_3  (
            .in0(N__10673),
            .in1(N__11354),
            .in2(N__10619),
            .in3(N__10918),
            .lcout(\uu2.w_addr_user_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNI24622_0_LC_8_5_4 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNI24622_0_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNI24622_0_LC_8_5_4 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \Lab_UT.dspStr.cnt_RNI24622_0_LC_8_5_4  (
            .in0(N__10920),
            .in1(N__8729),
            .in2(_gnd_net_),
            .in3(N__10143),
            .lcout(\Lab_UT.dspStr.cnt11_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dek.det_N_5_LC_8_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dek.det_N_5_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrluu0.dek.det_N_5_LC_8_5_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrluu0.dek.det_N_5_LC_8_5_5  (
            .in0(N__11983),
            .in1(N__11356),
            .in2(N__11420),
            .in3(N__11387),
            .lcout(),
            .ltout(\Lab_UT.dictrluu0.dek.det_NZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dek.det_N_LC_8_5_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dek.det_N_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrluu0.dek.det_N_LC_8_5_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrluu0.dek.det_N_LC_8_5_6  (
            .in0(N__11906),
            .in1(N__8936),
            .in2(N__8744),
            .in3(N__11457),
            .lcout(\Lab_UT.dicSelectLEDdisp ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_8_5_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_8_5_7 .LUT_INIT=16'b1110000011110101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_45_LC_8_5_7  (
            .in0(N__10674),
            .in1(N__11355),
            .in2(N__10620),
            .in3(N__10919),
            .lcout(\uu2.mem0.N_1476_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un27_m3_0_LC_8_6_0 .C_ON=1'b0;
    defparam \uu2.un27_m3_0_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un27_m3_0_LC_8_6_0 .LUT_INIT=16'b0001111100001010;
    LogicCell40 \uu2.un27_m3_0_LC_8_6_0  (
            .in0(N__10665),
            .in1(N__11357),
            .in2(N__10613),
            .in3(N__10917),
            .lcout(\uu2.un27_N_6_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNI11B71_3_LC_8_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNI11B71_3_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNI11B71_3_LC_8_6_1 .LUT_INIT=16'b0000000000110001;
    LogicCell40 \Lab_UT.dspStr.cnt_RNI11B71_3_LC_8_6_1  (
            .in0(N__13121),
            .in1(N__10595),
            .in2(N__11756),
            .in3(N__10666),
            .lcout(\Lab_UT.dspStr.cnt11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_m5_i_a3_2_LC_8_6_2 .C_ON=1'b0;
    defparam \uu2.w_m5_i_a3_2_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_m5_i_a3_2_LC_8_6_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.w_m5_i_a3_2_LC_8_6_2  (
            .in0(N__11455),
            .in1(N__11386),
            .in2(_gnd_net_),
            .in3(N__9053),
            .lcout(\uu2.w_m5_i_a3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrluu0.dek.det_N_4_LC_8_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrluu0.dek.det_N_4_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrluu0.dek.det_N_4_LC_8_6_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrluu0.dek.det_N_4_LC_8_6_3  (
            .in0(N__11330),
            .in1(N__10769),
            .in2(_gnd_net_),
            .in3(N__11944),
            .lcout(\Lab_UT.dictrluu0.dek.det_NZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_0_0_0_LC_8_6_4 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_0_0_0_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_0_0_0_LC_8_6_4 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \uu2.un1_w_user_lf_0_0_0_LC_8_6_4  (
            .in0(N__11456),
            .in1(N__10916),
            .in2(_gnd_net_),
            .in3(N__11329),
            .lcout(),
            .ltout(\uu2.un1_w_user_lf_0_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_0_LC_8_6_5 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_0_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_0_LC_8_6_5 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \uu2.un1_w_user_lf_0_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__10591),
            .in2(N__8930),
            .in3(N__10664),
            .lcout(\uu2.un1_w_user_lf_2 ),
            .ltout(\uu2.un1_w_user_lf_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNILDNK6_4_LC_8_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNILDNK6_4_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNILDNK6_4_LC_8_6_6 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \uu2.w_addr_user_RNILDNK6_4_LC_8_6_6  (
            .in0(N__8917),
            .in1(N__8803),
            .in2(N__8903),
            .in3(N__8900),
            .lcout(),
            .ltout(\uu2.w_addr_user_RNILDNK6Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIOM3NG_4_LC_8_6_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIOM3NG_4_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIOM3NG_4_LC_8_6_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \uu2.w_addr_user_RNIOM3NG_4_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__8893),
            .in2(N__8858),
            .in3(N__9017),
            .lcout(\uu2.un27_w_addr_user_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_5_a0_5_LC_8_7_0 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_5_a0_5_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_5_a0_5_LC_8_7_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uu2.un1_w_user_lf_5_a0_5_LC_8_7_0  (
            .in0(N__9052),
            .in1(N__8982),
            .in2(N__9008),
            .in3(N__11382),
            .lcout(),
            .ltout(\uu2.un1_w_user_lf_5_a0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_5_a0_LC_8_7_1 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_5_a0_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_5_a0_LC_8_7_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \uu2.un1_w_user_lf_5_a0_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__11409),
            .in2(N__8810),
            .in3(N__11882),
            .lcout(\uu2.un1_w_user_lf_5_aZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_1_rep1_LC_8_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_1_rep1_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_1_rep1_LC_8_7_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.dspStr.cnt_1_rep1_LC_8_7_2  (
            .in0(N__11054),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(Lab_UT_dspStr_cnt_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13418),
            .ce(),
            .sr(N__12303));
    defparam \Lab_UT.dspStr.cnt_2_rep1_LC_8_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_2_rep1_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_2_rep1_LC_8_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dspStr.cnt_2_rep1_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11513),
            .lcout(Lab_UT_dspStr_cnt_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13418),
            .ce(),
            .sr(N__12303));
    defparam \Lab_UT.dspStr.cnt_3_rep1_LC_8_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_3_rep1_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_3_rep1_LC_8_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dspStr.cnt_3_rep1_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11306),
            .lcout(Lab_UT_dspStr_cnt_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13418),
            .ce(),
            .sr(N__12303));
    defparam \Lab_UT.dspStr.cnt_3_rep1_RNIIV651_LC_8_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_3_rep1_RNIIV651_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_3_rep1_RNIIV651_LC_8_7_5 .LUT_INIT=16'b1011111111001100;
    LogicCell40 \Lab_UT.dspStr.cnt_3_rep1_RNIIV651_LC_8_7_5  (
            .in0(N__8981),
            .in1(N__8999),
            .in2(N__11323),
            .in3(N__9050),
            .lcout(Lab_UT_L3_tx_data_0_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_3_rep1_RNI05SQ_LC_8_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_3_rep1_RNI05SQ_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_3_rep1_RNI05SQ_LC_8_7_6 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \Lab_UT.dspStr.cnt_3_rep1_RNI05SQ_LC_8_7_6  (
            .in0(N__9051),
            .in1(_gnd_net_),
            .in2(N__9007),
            .in3(N__8980),
            .lcout(Lab_UT_dspStr_un36_dOut),
            .ltout(Lab_UT_dspStr_un36_dOut_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_1_LC_8_7_7 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_1_LC_8_7_7 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \uu2.un1_w_user_cr_1_LC_8_7_7  (
            .in0(N__11967),
            .in1(N__10963),
            .in2(N__9023),
            .in3(N__11023),
            .lcout(\uu2.un1_w_user_crZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un4_w_user_data_rdy_0_LC_8_8_0 .C_ON=1'b0;
    defparam \uu2.un4_w_user_data_rdy_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un4_w_user_data_rdy_0_LC_8_8_0 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \uu2.un4_w_user_data_rdy_0_LC_8_8_0  (
            .in0(N__9292),
            .in1(N__11088),
            .in2(N__8959),
            .in3(N__9313),
            .lcout(\uu2.un4_w_user_data_rdyZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un27_m3_LC_8_8_1 .C_ON=1'b0;
    defparam \uu2.un27_m3_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un27_m3_LC_8_8_1 .LUT_INIT=16'b0000001101110011;
    LogicCell40 \uu2.un27_m3_LC_8_8_1  (
            .in0(N__11448),
            .in1(N__10925),
            .in2(N__10618),
            .in3(N__8983),
            .lcout(),
            .ltout(\uu2.un27_N_6_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un27_w_addr_user_i_1_LC_8_8_2 .C_ON=1'b0;
    defparam \uu2.un27_w_addr_user_i_1_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.un27_w_addr_user_i_1_LC_8_8_2 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \uu2.un27_w_addr_user_i_1_LC_8_8_2  (
            .in0(N__9290),
            .in1(N__11086),
            .in2(N__9020),
            .in3(N__9311),
            .lcout(\uu2.un27_w_addr_user_iZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_3_rep1_RNIEPV31_LC_8_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_3_rep1_RNIEPV31_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_3_rep1_RNIEPV31_LC_8_8_3 .LUT_INIT=16'b1110111010100010;
    LogicCell40 \Lab_UT.dspStr.cnt_3_rep1_RNIEPV31_LC_8_8_3  (
            .in0(N__10935),
            .in1(N__9006),
            .in2(N__11458),
            .in3(N__8984),
            .lcout(L3_tx_data_0),
            .ltout(L3_tx_data_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIQKOV8_8_LC_8_8_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIQKOV8_8_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIQKOV8_8_LC_8_8_4 .LUT_INIT=16'b1111111111010101;
    LogicCell40 \uu2.w_addr_displaying_RNIQKOV8_8_LC_8_8_4  (
            .in0(N__9291),
            .in1(N__11087),
            .in2(N__9323),
            .in3(N__9899),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_RNIQKOV8Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIB9CMF_8_LC_8_8_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIB9CMF_8_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIB9CMF_8_LC_8_8_5 .LUT_INIT=16'b1110010011110101;
    LogicCell40 \uu2.w_addr_displaying_RNIB9CMF_8_LC_8_8_5  (
            .in0(N__9312),
            .in1(N__9902),
            .in2(N__9296),
            .in3(N__9293),
            .lcout(\uu2.un21_w_addr_displaying_i ),
            .ltout(\uu2.un21_w_addr_displaying_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_6_LC_8_8_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_6_LC_8_8_6 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_fast_6_LC_8_8_6 .LUT_INIT=16'b1101111111100000;
    LogicCell40 \uu2.w_addr_displaying_fast_6_LC_8_8_6  (
            .in0(N__11817),
            .in1(N__9900),
            .in2(N__9260),
            .in3(N__12098),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_6C_net ),
            .ce(),
            .sr(N__12283));
    defparam \uu2.mem0.ram512X8_inst_RNO_69_LC_8_9_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_69_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_69_LC_8_9_0 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_69_LC_8_9_0  (
            .in0(N__12871),
            .in1(N__13055),
            .in2(N__12998),
            .in3(N__13226),
            .lcout(\uu2.mem0.g0_i_a11_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_8_9_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_8_9_1 .LUT_INIT=16'b0101000000100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_55_LC_8_9_1  (
            .in0(N__13228),
            .in1(N__12991),
            .in2(N__13066),
            .in3(N__12874),
            .lcout(),
            .ltout(\uu2.mem0.g3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_8_9_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_8_9_2 .LUT_INIT=16'b1101010100000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_33_LC_8_9_2  (
            .in0(N__12086),
            .in1(N__9238),
            .in2(N__9167),
            .in3(N__9156),
            .lcout(\uu2.mem0.un1_segment4_0_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_70_LC_8_9_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_70_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_70_LC_8_9_3 .LUT_INIT=16'b0000100010000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_70_LC_8_9_3  (
            .in0(N__13225),
            .in1(N__12984),
            .in2(N__13065),
            .in3(N__12872),
            .lcout(\uu2.mem0.g0_i_a11_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_68_LC_8_9_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_68_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_68_LC_8_9_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_68_LC_8_9_4  (
            .in0(N__12873),
            .in1(_gnd_net_),
            .in2(N__12999),
            .in3(N__13227),
            .lcout(),
            .ltout(\uu2.mem0.g0_i_a11_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_8_9_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_8_9_5 .LUT_INIT=16'b0101011111111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_57_LC_8_9_5  (
            .in0(N__9616),
            .in1(N__11522),
            .in2(N__9065),
            .in3(N__9796),
            .lcout(\uu2.mem0.g0_i_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_0_LC_8_9_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_0_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_0_LC_8_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_fast_0_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__9617),
            .in2(_gnd_net_),
            .in3(N__12466),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_0C_net ),
            .ce(),
            .sr(N__12287));
    defparam \uu2.w_addr_displaying_fast_RNI3A1N_0_LC_8_9_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI3A1N_0_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI3A1N_0_LC_8_9_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI3A1N_0_LC_8_9_7  (
            .in0(N__9615),
            .in1(N__9409),
            .in2(N__11637),
            .in3(N__9338),
            .lcout(\uu2.Z_decfrac106_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_61_LC_8_10_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_61_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_61_LC_8_10_0 .LUT_INIT=16'b0010100000010100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_61_LC_8_10_0  (
            .in0(N__11627),
            .in1(N__9787),
            .in2(N__12357),
            .in3(N__10006),
            .lcout(\uu2.mem0.bitmap_pmux_1_1_i_a5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_63_LC_8_10_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_63_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_63_LC_8_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_63_LC_8_10_1  (
            .in0(N__9597),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9538),
            .lcout(),
            .ltout(\uu2.mem0.g1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_8_10_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_8_10_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_43_LC_8_10_2  (
            .in0(N__9428),
            .in1(N__9476),
            .in2(N__9470),
            .in3(N__9462),
            .lcout(\uu2.mem0.g0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_62_LC_8_10_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_62_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_62_LC_8_10_3 .LUT_INIT=16'b0010100000010100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_62_LC_8_10_3  (
            .in0(N__10005),
            .in1(N__9411),
            .in2(N__9344),
            .in3(N__11628),
            .lcout(\uu2.mem0.bitmap_pmux_1_1_i_a5_2_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIFM1N_1_LC_8_10_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIFM1N_1_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIFM1N_1_LC_8_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIFM1N_1_LC_8_10_4  (
            .in0(N__9412),
            .in1(N__9788),
            .in2(N__12358),
            .in3(N__9342),
            .lcout(\uu2.Z_decfrac105_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_1_LC_8_10_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_1_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_1_LC_8_10_5 .LUT_INIT=16'b0110101001101010;
    LogicCell40 \uu2.w_addr_displaying_fast_1_LC_8_10_5  (
            .in0(N__9343),
            .in1(N__12563),
            .in2(N__12508),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_1C_net ),
            .ce(),
            .sr(N__12289));
    defparam \uu2.w_addr_displaying_fast_3_LC_8_10_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_3_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_3_LC_8_10_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \uu2.w_addr_displaying_fast_3_LC_8_10_6  (
            .in0(N__11531),
            .in1(_gnd_net_),
            .in2(N__11638),
            .in3(N__12489),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_1C_net ),
            .ce(),
            .sr(N__12289));
    defparam \uu2.mem0.ram512X8_inst_RNO_65_LC_8_10_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_65_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_65_LC_8_10_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_65_LC_8_10_7  (
            .in0(N__10007),
            .in1(N__11629),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.mem0.Z_decfrac105_7_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_8_LC_8_11_1 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_8_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_8_LC_8_11_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_8_LC_8_11_1  (
            .in0(N__12773),
            .in1(N__9671),
            .in2(N__9761),
            .in3(N__9944),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_4_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_8_LC_8_11_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_LC_8_11_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uu2.w_addr_displaying_8_LC_8_11_2  (
            .in0(N__9945),
            .in1(_gnd_net_),
            .in2(N__9971),
            .in3(N__12486),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8C_net ),
            .ce(),
            .sr(N__12290));
    defparam \uu2.w_addr_displaying_RNI4K2N2_8_LC_8_11_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI4K2N2_8_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI4K2N2_8_LC_8_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI4K2N2_8_LC_8_11_3  (
            .in0(N__12769),
            .in1(N__9669),
            .in2(N__9760),
            .in3(N__9943),
            .lcout(\uu2.un15_w_data_displaying ),
            .ltout(\uu2.un15_w_data_displaying_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_6_LC_8_11_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_LC_8_11_4 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_6_LC_8_11_4 .LUT_INIT=16'b1111011011001100;
    LogicCell40 \uu2.w_addr_displaying_6_LC_8_11_4  (
            .in0(N__11818),
            .in1(N__9842),
            .in2(N__9875),
            .in3(N__12487),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8C_net ),
            .ce(),
            .sr(N__12290));
    defparam \uu2.w_addr_displaying_7_LC_8_11_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_LC_8_11_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_7_LC_8_11_5  (
            .in0(N__12485),
            .in1(N__9750),
            .in2(N__12797),
            .in3(N__9672),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8C_net ),
            .ce(),
            .sr(N__12290));
    defparam \uu2.w_addr_displaying_fast_7_LC_8_11_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_7_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_7_LC_8_11_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_displaying_fast_7_LC_8_11_6  (
            .in0(N__12787),
            .in1(N__9795),
            .in2(N__9762),
            .in3(N__12488),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8C_net ),
            .ce(),
            .sr(N__12290));
    defparam \uu2.vbuf_w_addr_displaying.result_1_fast_8_LC_8_11_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_fast_8_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_fast_8_LC_8_11_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_fast_8_LC_8_11_7  (
            .in0(N__12355),
            .in1(N__9749),
            .in2(N__12796),
            .in3(N__9670),
            .lcout(\uu2.w_addr_displaying_4_fast_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_0_LC_8_12_0 .C_ON=1'b1;
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_0_LC_8_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_RNO_0_0_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__13223),
            .in2(N__11729),
            .in3(N__11730),
            .lcout(\Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\Lab_UT.didpuu0.didpsones.un1_q_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_1_LC_8_12_1 .C_ON=1'b1;
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_1_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_1_LC_8_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_RNO_0_1_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__12867),
            .in2(_gnd_net_),
            .in3(N__10127),
            .lcout(\Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\Lab_UT.didpuu0.didpsones.un1_q_cry_0 ),
            .carryout(\Lab_UT.didpuu0.didpsones.un1_q_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_2_LC_8_12_2 .C_ON=1'b1;
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_2_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_2_LC_8_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_RNO_0_2_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__13040),
            .in2(_gnd_net_),
            .in3(N__10118),
            .lcout(\Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\Lab_UT.didpuu0.didpsones.un1_q_cry_1 ),
            .carryout(\Lab_UT.didpuu0.didpsones.un1_q_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_3_LC_8_12_3 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.didpsones.q_RNO_0_3_LC_8_12_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_RNO_0_3_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__12979),
            .in2(_gnd_net_),
            .in3(N__10115),
            .lcout(),
            .ltout(\Lab_UT.didpuu0.didpsones.q_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_3_LC_8_12_4 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_3_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpsones.q_3_LC_8_12_4 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_3_LC_8_12_4  (
            .in0(N__10079),
            .in1(N__10095),
            .in2(N__10112),
            .in3(N__11731),
            .lcout(Lab_UT_di_Sones_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13391),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_0_LC_8_12_5 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_0_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpsones.q_0_LC_8_12_5 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_0_LC_8_12_5  (
            .in0(N__10109),
            .in1(N__11719),
            .in2(N__10096),
            .in3(N__10077),
            .lcout(Lab_UT_di_Sones_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13391),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_2_LC_8_12_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_2_LC_8_12_6 .LUT_INIT=16'b0000101010101010;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_8_12_6  (
            .in0(N__10532),
            .in1(_gnd_net_),
            .in2(N__10284),
            .in3(N__10505),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13391),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.didpsones.q_1_LC_8_12_7 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.didpsones.q_1_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didpuu0.didpsones.q_1_LC_8_12_7 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \Lab_UT.didpuu0.didpsones.q_1_LC_8_12_7  (
            .in0(N__10103),
            .in1(N__11720),
            .in2(N__10097),
            .in3(N__10078),
            .lcout(Lab_UT_di_Sones_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13391),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_LC_8_13_0 .C_ON=1'b1;
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.un1_bitcount_cry_0_c_LC_8_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.un1_bitcount_cry_0_c_LC_8_13_0  (
            .in0(_gnd_net_),
            .in1(N__10034),
            .in2(N__10373),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\buart.Z_tx.un1_bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_1_LC_8_13_1 .C_ON=1'b1;
    defparam \buart.Z_tx.bitcount_RNO_0_1_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_1_LC_8_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_1_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__10331),
            .in2(N__10352),
            .in3(N__10022),
            .lcout(\buart.Z_tx.bitcount_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\buart.Z_tx.un1_bitcount_cry_0 ),
            .carryout(\buart.Z_tx.un1_bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_8_13_2 .C_ON=1'b1;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_8_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__10400),
            .in2(N__10394),
            .in3(N__10526),
            .lcout(\buart.Z_tx.bitcount_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.un1_bitcount_cry_1 ),
            .carryout(\buart.Z_tx.un1_bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_3_LC_8_13_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.bitcount_3_LC_8_13_3 .LUT_INIT=16'b1011001111101100;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_8_13_3  (
            .in0(N__10244),
            .in1(N__10178),
            .in2(N__10523),
            .in3(N__10403),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13387),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIM5O32_2_LC_8_13_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIM5O32_2_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIM5O32_2_LC_8_13_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIM5O32_2_LC_8_13_4  (
            .in0(N__10393),
            .in1(N__10240),
            .in2(_gnd_net_),
            .in3(N__10321),
            .lcout(\buart.Z_tx.bitcount_RNIM5O32Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_8_13_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIQOQA1_3_LC_8_13_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_tx.bitcount_RNIQOQA1_3_LC_8_13_5  (
            .in0(N__10389),
            .in1(N__10347),
            .in2(N__10193),
            .in3(N__10367),
            .lcout(buart__tx_uart_busy_0),
            .ltout(buart__tx_uart_busy_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIL4O32_1_LC_8_13_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIL4O32_1_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIL4O32_1_LC_8_13_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIL4O32_1_LC_8_13_6  (
            .in0(N__10348),
            .in1(_gnd_net_),
            .in2(N__10334),
            .in3(N__10320),
            .lcout(\buart.Z_tx.bitcount_RNIL4O32Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_8_13_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_8_13_7 .LUT_INIT=16'b1111010100001010;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_8_13_7  (
            .in0(N__10322),
            .in1(_gnd_net_),
            .in2(N__10274),
            .in3(N__10192),
            .lcout(\buart.Z_tx.un1_bitcount_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.secuu0.sec_clkD_LC_9_4_6 .C_ON=1'b0;
    defparam \Lab_UT.secuu0.sec_clkD_LC_9_4_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.secuu0.sec_clkD_LC_9_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.secuu0.sec_clkD_LC_9_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13117),
            .lcout(\Lab_UT.sec_clkD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13433),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_0_LC_9_5_0 .C_ON=1'b1;
    defparam \Lab_UT.dspStr.cnt_0_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_0_LC_9_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.dspStr.cnt_0_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__10144),
            .in2(N__10172),
            .in3(N__10168),
            .lcout(\Lab_UT.dspStr.cntZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\Lab_UT.dspStr.un1_cnt_3_cry_0 ),
            .clk(N__13431),
            .ce(),
            .sr(N__12306));
    defparam \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87E_LC_9_5_1 .C_ON=1'b1;
    defparam \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87E_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87E_LC_9_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87E_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__10924),
            .in2(_gnd_net_),
            .in3(N__10952),
            .lcout(\Lab_UT.dspStr.un1_cnt_3_cry_0_c_RNIS87EZ0 ),
            .ltout(),
            .carryin(\Lab_UT.dspStr.un1_cnt_3_cry_0 ),
            .carryout(\Lab_UT.dspStr.un1_cnt_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8E_LC_9_5_2 .C_ON=1'b1;
    defparam \Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8E_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8E_LC_9_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8E_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__10679),
            .in2(_gnd_net_),
            .in3(N__10949),
            .lcout(\Lab_UT.dspStr.un1_cnt_3_cry_1_c_RNIUB8EZ0 ),
            .ltout(),
            .carryin(\Lab_UT.dspStr.un1_cnt_3_cry_1 ),
            .carryout(\Lab_UT.dspStr.un1_cnt_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9E_LC_9_5_3 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9E_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9E_LC_9_5_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9E_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__10579),
            .in2(_gnd_net_),
            .in3(N__10946),
            .lcout(\Lab_UT.dspStr.un1_cnt_3_cry_2_c_RNI0F9EZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_1_LC_9_5_4 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_1_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_1_LC_9_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dspStr.cnt_1_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11046),
            .lcout(Lab_UT_dspStr_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13431),
            .ce(),
            .sr(N__12306));
    defparam \Lab_UT.Lab3U01.q_0_LC_9_6_0 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U01.q_0_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U01.q_0_LC_9_6_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.Lab3U01.q_0_LC_9_6_0  (
            .in0(N__10763),
            .in1(N__10874),
            .in2(N__10829),
            .in3(N__10790),
            .lcout(\Lab_UT.rx_data_rdy ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13428),
            .ce(),
            .sr(N__12305));
    defparam \resetGen.un3_reset_count_i_a3_4_LC_9_6_1 .C_ON=1'b0;
    defparam \resetGen.un3_reset_count_i_a3_4_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \resetGen.un3_reset_count_i_a3_4_LC_9_6_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \resetGen.un3_reset_count_i_a3_4_LC_9_6_1  (
            .in0(N__13511),
            .in1(N__13486),
            .in2(_gnd_net_),
            .in3(N__10762),
            .lcout(\resetGen.un3_reset_count_i_a3Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_RNIN6202_3_LC_9_6_2 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_RNIN6202_3_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_RNIN6202_3_LC_9_6_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \Lab_UT.dspStr.cnt_RNIN6202_3_LC_9_6_2  (
            .in0(N__10578),
            .in1(N__10675),
            .in2(_gnd_net_),
            .in3(N__11114),
            .lcout(Lab_UT_L3_tx_data_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_2_LC_9_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_2_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_2_LC_9_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dspStr.cnt_2_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11502),
            .lcout(Lab_UT_dspStr_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13428),
            .ce(),
            .sr(N__12305));
    defparam \Lab_UT.dspStr.cnt_3_LC_9_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_3_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_3_LC_9_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.dspStr.cnt_3_LC_9_6_4  (
            .in0(N__11298),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(Lab_UT_dspStr_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13428),
            .ce(),
            .sr(N__12305));
    defparam \Lab_UT.dspStr.cnt_fast_3_LC_9_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_fast_3_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_fast_3_LC_9_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dspStr.cnt_fast_3_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11299),
            .lcout(\Lab_UT.dspStr.cnt_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13428),
            .ce(),
            .sr(N__12305));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_9_6_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_9_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_9_6_7  (
            .in0(N__11285),
            .in1(N__12584),
            .in2(_gnd_net_),
            .in3(N__11213),
            .lcout(\uu2.mem0.w_addr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_fast_RNIU9551_1_LC_9_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_fast_RNIU9551_1_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_fast_RNIU9551_1_LC_9_7_0 .LUT_INIT=16'b1111001001011111;
    LogicCell40 \Lab_UT.dspStr.cnt_fast_RNIU9551_1_LC_9_7_0  (
            .in0(N__11008),
            .in1(N__11934),
            .in2(N__11489),
            .in3(N__10987),
            .lcout(),
            .ltout(Lab_UT_L3_tx_data_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_4_LC_9_7_1 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_4_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_4_LC_9_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.un1_w_user_cr_4_LC_9_7_1  (
            .in0(N__11066),
            .in1(N__11060),
            .in2(N__11117),
            .in3(N__11113),
            .lcout(\uu2.un1_w_user_crZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_fast_RNIQ5551_1_LC_9_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_fast_RNIQ5551_1_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_fast_RNIQ5551_1_LC_9_7_2 .LUT_INIT=16'b1111011110101111;
    LogicCell40 \Lab_UT.dspStr.cnt_fast_RNIQ5551_1_LC_9_7_2  (
            .in0(N__11007),
            .in1(N__11408),
            .in2(N__11488),
            .in3(N__10986),
            .lcout(Lab_UT_L3_tx_data_0_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_fast_RNIS7551_1_LC_9_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_fast_RNIS7551_1_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_fast_RNIS7551_1_LC_9_7_3 .LUT_INIT=16'b1111001110110011;
    LogicCell40 \Lab_UT.dspStr.cnt_fast_RNIS7551_1_LC_9_7_3  (
            .in0(N__11343),
            .in1(N__11005),
            .in2(N__10988),
            .in3(N__11476),
            .lcout(Lab_UT_L3_tx_data_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_fast_1_LC_9_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_fast_1_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_fast_1_LC_9_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dspStr.cnt_fast_1_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11053),
            .lcout(\Lab_UT.dspStr.cnt_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13425),
            .ce(),
            .sr(N__12304));
    defparam \Lab_UT.dspStr.cnt_fast_RNIR6551_1_LC_9_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_fast_RNIR6551_1_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_fast_RNIR6551_1_LC_9_7_5 .LUT_INIT=16'b1010101010000101;
    LogicCell40 \Lab_UT.dspStr.cnt_fast_RNIR6551_1_LC_9_7_5  (
            .in0(N__10984),
            .in1(N__11378),
            .in2(N__11012),
            .in3(N__11483),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_fast_RNIT8551_1_LC_9_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_fast_RNIT8551_1_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dspStr.cnt_fast_RNIT8551_1_LC_9_7_6 .LUT_INIT=16'b1101001111011011;
    LogicCell40 \Lab_UT.dspStr.cnt_fast_RNIT8551_1_LC_9_7_6  (
            .in0(N__11006),
            .in1(N__10985),
            .in2(N__11487),
            .in3(N__11898),
            .lcout(Lab_UT_L3_tx_data_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dspStr.cnt_fast_2_LC_9_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dspStr.cnt_fast_2_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dspStr.cnt_fast_2_LC_9_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dspStr.cnt_fast_2_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11509),
            .lcout(\Lab_UT.dspStr.cnt_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13425),
            .ce(),
            .sr(N__12304));
    defparam \Lab_UT.Lab3U00.q_esr_0_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_0_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_0_LC_9_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_0_LC_9_8_0  (
            .in0(N__12206),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(Lab_UT_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(N__11765),
            .sr(N__12300));
    defparam \Lab_UT.Lab3U00.q_esr_1_LC_9_8_1 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_1_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_1_LC_9_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_1_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12191),
            .lcout(Lab_UT_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(N__11765),
            .sr(N__12300));
    defparam \Lab_UT.Lab3U00.q_esr_2_LC_9_8_2 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_2_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_2_LC_9_8_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_2_LC_9_8_2  (
            .in0(N__13462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(Lab_UT_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(N__11765),
            .sr(N__12300));
    defparam \Lab_UT.Lab3U00.q_esr_3_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_3_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_3_LC_9_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_3_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13487),
            .lcout(Lab_UT_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(N__11765),
            .sr(N__12300));
    defparam \Lab_UT.Lab3U00.q_esr_4_LC_9_8_4 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_4_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_4_LC_9_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_4_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13510),
            .lcout(Lab_UT_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(N__11765),
            .sr(N__12300));
    defparam \Lab_UT.Lab3U00.q_esr_5_LC_9_8_5 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_5_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_5_LC_9_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_5_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12116),
            .lcout(Lab_UT_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(N__11765),
            .sr(N__12300));
    defparam \Lab_UT.Lab3U00.q_esr_6_LC_9_8_6 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_6_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_6_LC_9_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_6_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12137),
            .lcout(Lab_UT_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(N__11765),
            .sr(N__12300));
    defparam \Lab_UT.Lab3U00.q_esr_7_LC_9_8_7 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_7_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.Lab3U00.q_esr_7_LC_9_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_7_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12173),
            .lcout(Lab_UT_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13419),
            .ce(N__11765),
            .sr(N__12300));
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_9_9_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_9_9_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_54_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__12097),
            .in2(_gnd_net_),
            .in3(N__12613),
            .lcout(\uu2.mem0.N_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_3_LC_9_9_1 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_3_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_3_LC_9_9_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_3_LC_9_9_1  (
            .in0(N__11590),
            .in1(N__11695),
            .in2(N__12585),
            .in3(N__12080),
            .lcout(\uu2.w_addr_displaying_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_5_a0_4_LC_9_9_2 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_5_a0_4_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_5_a0_4_LC_9_9_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uu2.un1_w_user_lf_5_a0_4_LC_9_9_2  (
            .in0(N__11966),
            .in1(N__11924),
            .in2(_gnd_net_),
            .in3(N__11899),
            .lcout(\uu2.un1_w_user_lf_5_a0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_6__un437_ci_LC_9_9_3 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_6__un437_ci_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_6__un437_ci_LC_9_9_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.vbuf_w_addr_displaying.counter_gen_label_6__un437_ci_LC_9_9_3  (
            .in0(N__12804),
            .in1(N__11873),
            .in2(_gnd_net_),
            .in3(N__12706),
            .lcout(\uu2.un437_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.Lab3U00.q_esr_ctle_7_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.Lab3U00.q_esr_ctle_7_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.Lab3U00.q_esr_ctle_7_LC_9_9_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Lab_UT.Lab3U00.q_esr_ctle_7_LC_9_9_4  (
            .in0(N__11795),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12323),
            .lcout(\Lab_UT.Lab3U00.bu_rx_data_rdy_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.clkSecStrb_LC_9_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.clkSecStrb_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.clkSecStrb_LC_9_9_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.didpuu0.clkSecStrb_LC_9_9_5  (
            .in0(N__13136),
            .in1(N__11755),
            .in2(_gnd_net_),
            .in3(N__13168),
            .lcout(\Lab_UT.didpuu0.clkSecStrbZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_fast_3_LC_9_9_6 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_fast_3_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_fast_3_LC_9_9_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_fast_3_LC_9_9_6  (
            .in0(N__11696),
            .in1(N__12561),
            .in2(N__11639),
            .in3(N__11591),
            .lcout(\uu2.w_addr_displaying_4_fast_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_67_LC_9_9_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_67_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_67_LC_9_9_7 .LUT_INIT=16'b0000001010101000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_67_LC_9_9_7  (
            .in0(N__13054),
            .in1(N__12881),
            .in2(N__13000),
            .in3(N__13232),
            .lcout(\uu2.mem0.g0_i_a11_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_5_LC_9_10_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_5_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_5_LC_9_10_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_displaying_fast_5_LC_9_10_0  (
            .in0(N__12495),
            .in1(N__12614),
            .in2(N__12809),
            .in3(N__12710),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_5C_net ),
            .ce(),
            .sr(N__12291));
    defparam \uu2.w_addr_displaying_0_LC_9_10_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_9_10_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_0_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__12562),
            .in2(_gnd_net_),
            .in3(N__12496),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_5C_net ),
            .ce(),
            .sr(N__12291));
    defparam \uu2.w_addr_displaying_fast_8_LC_9_10_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_8_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_8_LC_9_10_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.w_addr_displaying_fast_8_LC_9_10_2  (
            .in0(N__12494),
            .in1(N__12377),
            .in2(_gnd_net_),
            .in3(N__12356),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_5C_net ),
            .ce(),
            .sr(N__12291));
    defparam \resetGen.un3_reset_count_i_a3_5_LC_9_11_0 .C_ON=1'b0;
    defparam \resetGen.un3_reset_count_i_a3_5_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \resetGen.un3_reset_count_i_a3_5_LC_9_11_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \resetGen.un3_reset_count_i_a3_5_LC_9_11_0  (
            .in0(N__12111),
            .in1(N__12186),
            .in2(N__12136),
            .in3(N__12202),
            .lcout(\resetGen.un3_reset_count_i_a3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_LC_9_11_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_0_LC_9_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_LC_9_11_1  (
            .in0(N__12187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13402),
            .ce(N__13259),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_LC_9_11_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_1_LC_9_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13452),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13402),
            .ce(N__13259),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_5_LC_9_11_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_5_LC_9_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12132),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13402),
            .ce(N__13259),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_6_LC_9_11_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_6_LC_9_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12168),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13402),
            .ce(N__13259),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_4_LC_9_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_4_LC_9_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_4_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12112),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13402),
            .ce(N__13259),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_3_LC_9_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_3_LC_9_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13506),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13402),
            .ce(N__13259),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_2_LC_9_11_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.shifter_2_LC_9_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13479),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13402),
            .ce(N__13259),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_0_LC_9_12_5 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_0_LC_9_12_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.L3_led_1_0_LC_9_12_5  (
            .in0(N__12919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13224),
            .lcout(led_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.o_oneSecPluse_LC_11_9_6 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.o_oneSecPluse_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.o_oneSecPluse_LC_11_9_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didpuu0.o_oneSecPluse_LC_11_9_6  (
            .in0(N__13169),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13144),
            .lcout(led_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_2_LC_11_11_2 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_2_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_2_LC_11_11_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.L3_led_1_2_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__12914),
            .in2(_gnd_net_),
            .in3(N__13067),
            .lcout(led_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_3_LC_11_11_3 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_3_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_3_LC_11_11_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.L3_led_1_3_LC_11_11_3  (
            .in0(N__12915),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13001),
            .lcout(led_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_1_LC_11_12_1 .C_ON=1'b0;
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_1_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didpuu0.ledDisp00.L3_led_1_1_LC_11_12_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.didpuu0.ledDisp00.L3_led_1_1_LC_11_12_1  (
            .in0(N__12923),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12880),
            .lcout(led_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // latticehx1k
